// Verilog netlist created by TD v5.0.27252
// Sat May 22 05:13:07 2021

`timescale 1ns / 1ps
module font_ram  // font_ram.v(14)
  (
  addra,
  clka,
  dia,
  wea,
  doa
  );

  input [14:0] addra;  // font_ram.v(29)
  input clka;  // font_ram.v(31)
  input [15:0] dia;  // font_ram.v(28)
  input wea;  // font_ram.v(30)
  output [15:0] doa;  // font_ram.v(26)

  parameter ADDR_WIDTH_A = 15;
  parameter ADDR_WIDTH_B = 15;
  parameter DATA_DEPTH_A = 20480;
  parameter DATA_DEPTH_B = 20480;
  parameter DATA_WIDTH_A = 16;
  parameter DATA_WIDTH_B = 16;
  parameter REGMODE_A = "NOREG";
  parameter WRITEMODE_A = "NORMAL";
  wire [0:2] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b0/B1_0 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b1/B1_0 ;
  wire  \inst_doa_mux_b10/B0_0 ;
  wire  \inst_doa_mux_b10/B0_1 ;
  wire  \inst_doa_mux_b10/B1_0 ;
  wire  \inst_doa_mux_b11/B0_0 ;
  wire  \inst_doa_mux_b11/B0_1 ;
  wire  \inst_doa_mux_b11/B1_0 ;
  wire  \inst_doa_mux_b12/B0_0 ;
  wire  \inst_doa_mux_b12/B0_1 ;
  wire  \inst_doa_mux_b12/B1_0 ;
  wire  \inst_doa_mux_b13/B0_0 ;
  wire  \inst_doa_mux_b13/B0_1 ;
  wire  \inst_doa_mux_b13/B1_0 ;
  wire  \inst_doa_mux_b14/B0_0 ;
  wire  \inst_doa_mux_b14/B0_1 ;
  wire  \inst_doa_mux_b14/B1_0 ;
  wire  \inst_doa_mux_b15/B0_0 ;
  wire  \inst_doa_mux_b15/B0_1 ;
  wire  \inst_doa_mux_b15/B1_0 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b2/B1_0 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b3/B1_0 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b4/B1_0 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b5/B1_0 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b6/B1_0 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire  \inst_doa_mux_b7/B1_0 ;
  wire  \inst_doa_mux_b8/B0_0 ;
  wire  \inst_doa_mux_b8/B0_1 ;
  wire  \inst_doa_mux_b8/B1_0 ;
  wire  \inst_doa_mux_b9/B0_0 ;
  wire  \inst_doa_mux_b9/B0_1 ;
  wire  \inst_doa_mux_b9/B1_0 ;
  wire \and_Naddra[12]_Naddr_o ;
  wire \and_Naddra[12]_Naddr_o_al_n16 ;
  wire \and_Naddra[12]_addra_o ;
  wire \and_addra[12]_Naddra_o ;
  wire \and_addra[12]_addra[_o ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i0_008;
  wire inst_doa_i0_009;
  wire inst_doa_i0_010;
  wire inst_doa_i0_011;
  wire inst_doa_i0_012;
  wire inst_doa_i0_013;
  wire inst_doa_i0_014;
  wire inst_doa_i0_015;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i1_008;
  wire inst_doa_i1_009;
  wire inst_doa_i1_010;
  wire inst_doa_i1_011;
  wire inst_doa_i1_012;
  wire inst_doa_i1_013;
  wire inst_doa_i1_014;
  wire inst_doa_i1_015;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;
  wire inst_doa_i2_008;
  wire inst_doa_i2_009;
  wire inst_doa_i2_010;
  wire inst_doa_i2_011;
  wire inst_doa_i2_012;
  wire inst_doa_i2_013;
  wire inst_doa_i2_014;
  wire inst_doa_i2_015;
  wire inst_doa_i3_000;
  wire inst_doa_i3_001;
  wire inst_doa_i3_002;
  wire inst_doa_i3_003;
  wire inst_doa_i3_004;
  wire inst_doa_i3_005;
  wire inst_doa_i3_006;
  wire inst_doa_i3_007;
  wire inst_doa_i3_008;
  wire inst_doa_i3_009;
  wire inst_doa_i3_010;
  wire inst_doa_i3_011;
  wire inst_doa_i3_012;
  wire inst_doa_i3_013;
  wire inst_doa_i3_014;
  wire inst_doa_i3_015;
  wire inst_doa_i4_000;
  wire inst_doa_i4_001;
  wire inst_doa_i4_002;
  wire inst_doa_i4_003;
  wire inst_doa_i4_004;
  wire inst_doa_i4_005;
  wire inst_doa_i4_006;
  wire inst_doa_i4_007;
  wire inst_doa_i4_008;
  wire inst_doa_i4_009;
  wire inst_doa_i4_010;
  wire inst_doa_i4_011;
  wire inst_doa_i4_012;
  wire inst_doa_i4_013;
  wire inst_doa_i4_014;
  wire inst_doa_i4_015;
  wire wea_neg;

  AL_DFF_X addra_pipe_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[12]),
    .en(wea_neg),
    .sr(1'b0),
    .ss(1'b0),
    .q(addra_piped[0]));
  AL_DFF_X addra_pipe_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[13]),
    .en(wea_neg),
    .sr(1'b0),
    .ss(1'b0),
    .q(addra_piped[1]));
  AL_DFF_X addra_pipe_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[14]),
    .en(wea_neg),
    .sr(1'b0),
    .ss(1'b0),
    .q(addra_piped[2]));
  and \and_Naddra[12]_Naddr  (\and_Naddra[12]_Naddr_o , ~addra[12], ~addra[13], ~addra[14]);
  and \and_Naddra[12]_Naddr_al_u16  (\and_Naddra[12]_Naddr_o_al_n16 , ~addra[12], ~addra[13], addra[14]);
  and \and_Naddra[12]_addra  (\and_Naddra[12]_addra_o , ~addra[12], addra[13], ~addra[14]);
  and \and_addra[12]_Naddra  (\and_addra[12]_Naddra_o , addra[12], ~addra[13], ~addra[14]);
  and \and_addra[12]_addra[  (\and_addra[12]_addra[_o , addra[12], addra[13], ~addra[14]);
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=16;working_depth=4096;working_width=8;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h404040800000000000000000001E101010100080404040400000000000000000),
    .INIT_01(256'h0000000000242418242400000000008000000000000000000012121E12120080),
    .INIT_02(256'h1038008040404080000000000000000000242418242400000000008000000000),
    .INIT_03(256'h0000000000000000000A1412120C004040C04040000000000000000000101010),
    .INIT_04(256'h001E1010101000C0000000C0000000000000000000121418141200C0000000C0),
    .INIT_05(256'h80808000000000000000000000000000E0106080700000000000000000000000),
    .INIT_06(256'h00000000000000008080C080F000000000000000000000000038243824380080),
    .INIT_07(256'h8080C080F0000000000000000000000000000000202020207000000000000000),
    .INIT_08(256'h00000000000000000000000090A0E090E0000000000000000000000000000000),
    .INIT_09(256'h00000000E0404040E0000000000000000000000000000000E010608070000000),
    .INIT_0A(256'h000000C00000000000000000001E1018101E00C0000000000000000000000000),
    .INIT_0B(256'h00000000001C1008041800C0000000C00000000000000000001C0808180800C0),
    .INIT_0C(256'h141400C0000000C0000000000000000000180408041800C0000000C000000000),
    .INIT_0D(256'h0000000000000000001214181412004040C0408000000000000000000004041C),
    .INIT_0E(256'h001C121C121C00000000008000000000000000000024242C3424000000008080),
    .INIT_0F(256'h880000000000000000000000001212161A12004040C040800000000000000000),
    .INIT_10(256'h00000000001C121C121C0080404040400000000000000000000000008888A8D8),
    .INIT_11(256'hE0106080700000000000000000000000000E1010100E0080408000C000000000),
    .INIT_12(256'h000000000000000000000000E010608070000000000000000000000000000000),
    .INIT_13(256'h00000000E010608070000000000000000000000000000000E010608070000000),
    .INIT_14(256'h0000008080808080800000000000000000000000000000000000000000000000),
    .INIT_15(256'hC0C00000000000000000000000000000C0C0C0C0C0C000000000000000000000),
    .INIT_16(256'hC0E070303070E0C0000030F0E000000000000000C0C0C0C0F0F0C0C0F0F0C0C0),
    .INIT_17(256'h00000000000000000000000060F0F06000000080C0E070300000000000000000),
    .INIT_18(256'h00000000000000000000000000000000000000000000000030F0E0E0F0300000),
    .INIT_19(256'hC0C0C0C0C0C0800000000000000000C0C08000000000000000000080C0C00000),
    .INIT_1A(256'h000000000000000000003070E0C08080C0E070300000000000000000000080C0),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000F0F000000000),
    .INIT_1C(256'h00000000000000000000000000000000F0F00000000000000000000000000000),
    .INIT_1D(256'h00000000000000000080C0E06070381C0C060703000000000000000000000000),
    .INIT_1E(256'h000000000000000000000000000000000080C0E0703030303070E0C080000000),
    .INIT_1F(256'hF0F0000000000000F0F000000000C0E070303070E0C000000000000000000000),
    .INIT_20(256'hC0C0C0C0F0F0C0C0C0C0C0C0C0C0000000000000C0E070303070E0C0C0E07030),
    .INIT_21(256'h00000000C0C0000000000000C0E0703030303070E0C00000F0F0000000000000),
    .INIT_22(256'h000000000000000000000080C0E07030F0F0000000000000C0E070303070E0C0),
    .INIT_23(256'h3030B0F070303070E0C0000000000000C0E070303070E0E070303070E0C00000),
    .INIT_24(256'h00000000000000000000000000000000000000000000000000000000C0E07030),
    .INIT_25(256'h70E0C080000000000080C0E07030000000000000000000000000000000000000),
    .INIT_26(256'h80000000000000000000000000000000F0F00000F0F000000000000000000030),
    .INIT_27(256'h00000000000000000080C0E070303070E0C00000000000000000000080C0E0C0),
    .INIT_28(256'hF0F0303030303070E0C0000000000000C0C00000E0F03030F0F03070E0C00000),
    .INIT_29(256'hE0C0000000000000C0E070303070E0E070303070E0C000000000000030303030),
    .INIT_2A(256'hC0E070303030303030303070E0C0000000000000C0E070300000000000003070),
    .INIT_2B(256'h00000000F0F0000000000000F0F000000000000000000000F0F0000000000000),
    .INIT_2C(256'h00000000E0F03030F0F0000000003070E0C00000000000000000000000000000),
    .INIT_2D(256'h0000000000000000C0C0000000000000303030303030F0F03030303030300000),
    .INIT_2E(256'h70300000000000000080C0C0C0C0C0C0C0C0C0C0F0F0000000000000C0C00000),
    .INIT_2F(256'hF0F00000000000000000000000000000000000003070E0C0800000000080C0E0),
    .INIT_30(256'h303030303030000000000000303030303030303030B0F0F07030000000000000),
    .INIT_31(256'h00000000C0E070303030303030303070E0C000000000000030303070F0F0B030),
    .INIT_32(256'hB030303030303070E0C0000000000000000000000000C0E070303070E0C00000),
    .INIT_33(256'hE0C00000000000003070E0C08000C0E070303070E0C00000000000003070E0C0),
    .INIT_34(256'h000000000000000000000000F0F0000000000000C0E070303070E0C000003070),
    .INIT_35(256'h703030303030000000000000C0E0703030303030303030303030000000000000),
    .INIT_36(256'h00000000C0E0F0303030303030303030303000000000000000008080C0C0C060),
    .INIT_37(256'h00008080C0E06070303000000000000030307060E0C08080C0E0607030300000),
    .INIT_38(256'hF0F0000000000000F0F0000000000080C0E07030F0F000000000000000000000),
    .INIT_39(256'h1C387060E0C080000000000000000000000000F0F00000000000000000000000),
    .INIT_3A(256'h3070E0C080000000000000C0C0C0C0C0C0C0C0C0C0C0C0C0C0C000000307060E),
    .INIT_3B(256'h0000FCFC00000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h7070F0F0B0300000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000C0E0703030303070E0C00000000000000000000030B0F0F0),
    .INIT_3E(256'hF0F0303030303030F0F030303030000000000000C0C0000000000000C0C00000),
    .INIT_3F(256'h00003070E0C0000000000000E0E00000F0F03070E0C000000000000000000000),
    .INIT_40(256'hC0E070303030F0F030303030F0F0000000000000000000000000000000000000),
    .INIT_41(256'h000000000000000000000000000000003030303030303070E0C0000000000000),
    .INIT_42(256'h000000000080C0C0C0C0C0C0C0C0C0C0C0C00000C0C0000000000000C0C00000),
    .INIT_43(256'hC0C00000000000000000000000000000000000003070E0C08080C0E070300000),
    .INIT_44(256'hE0C00000000000000000000030303030303030F0E0C000000000000000000000),
    .INIT_45(256'h00000000C0E0703030303070E0C0000000000000000000003030303030303070),
    .INIT_46(256'h30303030F0F000000000000000000000C0E0703030303070E0C0000000000000),
    .INIT_47(256'h00000000000000000000000000003070E0C000000000000030303030F0F03030),
    .INIT_48(256'hC0C0000000000000C0C000000000000000000000C0E07070E0C00000E0E00000),
    .INIT_49(256'h30300000000000000000000030B0F0F070303030303000000000000000000000),
    .INIT_4A(256'h00000000C0E0F03030303030303000000000000000000000008080C0C0E06070),
    .INIT_4B(256'hF0F070303030000000000000000000003070E0C08080C0E07030000000000000),
    .INIT_4C(256'hF0F0000000000000F0F000000080C0E0F0F0000000000000C0E07030303030B0),
    .INIT_4D(256'h00000000000000000000000000000000000000F0F08000000000000000000080),
    .INIT_4E(256'h00000000000000000000000080C0C0C0E0703870E0C0C0C08000000000000000),
    .INIT_4F(256'h0000000000000000000000C6C6C6D6FEEEC600000000000000000000F0F89C0C),
    .INIT_50(256'hE0E0E0B0301800000000000000000000000000000000000000003070E0C00000),
    .INIT_51(256'hE00000000000000080C0E06060E0C08080C0C0C080000000000000001830B0E0),
    .INIT_52(256'h0008D0E070303070E0D0080000000000000000000000000000000000006060E0),
    .INIT_53(256'h0000000000000000000000003070E0C0C0C0F0F0000000000000000000000000),
    .INIT_54(256'h00000000F0F030300000808000003030F0F00000000000000000000000000000),
    .INIT_55(256'h8080E0F0301800000000000000000000000000000000000000000000C0C00000),
    .INIT_56(256'hC08000000000000000000000000000E0F0381800000000000000000000000080),
    .INIT_57(256'hFCFC30B0F0F0703000000000000000000000000080C0E0603030F0F0303060E0),
    .INIT_58(256'h00000000000000000000FCFCC0E070381C9CF8F0000000000000000000003030),
    .INIT_59(256'h00000000F0F0C0C0E0703030303070E0C000000000003030FCFC30B0F0F07030),
    .INIT_5A(256'h6060C0C08080000000000000000000000080C0C0C0C0C080800000C0E0600000),
    .INIT_5B(256'h6000000000000000C0C00000C0C00000C0C000000000000000000000F8F83030),
    .INIT_5C(256'h00000000000000000000000080C0C0000000000080C0E0606060606060606060),
    .INIT_5D(256'h70000000000000000000000060606060606060606060E0C08000000000000000),
    .INIT_5E(256'h00000000000000000000000000000000000000000000000070F8DC8C8C8C9CF8),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h70E0C080000000000080C0E07030000000000000000000000000000000000000),
    .INIT_62(256'h80000000000000000000000000000000F0F00000E0F0381800000000C0C08030),
    .INIT_63(256'h000000000000000000000000000000000000000000000080C0E0703080C0E0C0),
    .INIT_64(256'hC0C0C08080800000808000000000000000000000000000000000000000000000),
    .INIT_65(256'hE0C000000000C0C0F0F0C0C0C0C0C0C0F0F0C0C0000000000000000080C0C0C0),
    .INIT_66(256'hC0E070308080000080803070E0C0000000000000F0F030300000C0C0000030F0),
    .INIT_67(256'hF0F0000080C0C00000000000C0808080F080C0C0607030381818000000000000),
    .INIT_68(256'h00000000C0E07070E0F03838F0E00000F0F0000000000000C0E07030F0F00000),
    .INIT_69(256'h06060606C6CE0C3CF8E0000000000000C0E07070E0C00000E0E0000080C0C000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000E0F83C0CCEC6),
    .INIT_6B(256'h1818181818F8F80000000000000000000000000000CCDCB870E070B8DCCC0000),
    .INIT_6C(256'hE6CE0C3CF8E0000000000000000000000000B0F0703070F0B000000000000000),
    .INIT_6D(256'h00000000000000000000000000000000C0C000000000E0F83C0C6E66C6C6E666),
    .INIT_6E(256'h00000000F0F0000000000000000000000000000000000080C0E060E0C0800000),
    .INIT_6F(256'hC080000000000000000000000000C0C0000080C0C080000000000000F0F00000),
    .INIT_70(256'hF0F030100080C0E0F0F0000080C0C0000000000000000000000080C0C08080C0),
    .INIT_71(256'hB0B0B0B0FCFC000000000000000080C0E0606060606000000000000000000000),
    .INIT_72(256'h0000000000000000008080000000000000000000000000B0B0B0B0B0B0B0B0B0),
    .INIT_73(256'h00000000000000000000000000000000F0F000000080C0E0F0F0000080C0C000),
    .INIT_74(256'h0000000000000000000000000000000080808080000000000000000000000000),
    .INIT_75(256'hF0F000000000C0C000000000F0F0000000000000000080C0E070E0C080000000),
    .INIT_76(256'h70300000C0C0000000000000F8F80000FCFC0C9CF8F000000000000000000000),
    .INIT_77(256'h00000000C0E0703000000000000000000000000000000000000000000080C0E0),
    .INIT_78(256'hF0303070E0C0000080C0C00000000000303030F0F0303070E0C0000000000000),
    .INIT_79(256'hC060600000000000303030F0F0303070E0C000C0C080000000000000303030F0),
    .INIT_7A(256'h303030F0F0303070E0C00000C0C0000000000000303030F0F0303070E0C00000),
    .INIT_7B(256'h80808080F8F8000000000000303030F0F0303070E0C000008080000000000000),
    .INIT_7C(256'h00000000C0E070300000000000003070E0C0000000000000F8F880808080E0E0),
    .INIT_7D(256'h00000000E0E0000080C0C00000000000E0E0000000000000E0E0000000000000),
    .INIT_7E(256'hC0C0000000000000E0E0000000000000E0E000C0C080000000000000E0E00000),
    .INIT_7F(256'hC0C0000000000000C0C000000000000000000000E0E0000000000000E0E00000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_20480x16_sub_000000_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_Naddra[12]_Naddr_o ),
    .dia({open_n51,open_n52,open_n53,open_n54,open_n55,open_n56,open_n57,open_n58,dia[7:0]}),
    .wea(wea),
    .doa({open_n80,open_n81,open_n82,open_n83,open_n84,open_n85,open_n86,open_n87,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}));
  // address_offset=0;data_offset=8;depth=4096;width=8;num_section=1;width_per_section=8;section_size=16;working_depth=4096;working_width=8;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0202020100700830403800000000000000000001020202020048485868480000),
    .INIT_01(256'h4078000000000000000000010101010300700830403800000000000000000001),
    .INIT_02(256'h0000000102020201007840604078000000000000000000010101010300784060),
    .INIT_03(256'h0048487848300000000000000000000202020302007840604078000000000000),
    .INIT_04(256'h0000000000000003020302030070487048700000000000000000000102020201),
    .INIT_05(256'h040704030020202020700000000000000000000000001C121C121C0000000000),
    .INIT_06(256'h00000000000000000000000000001E1010101000000000000000000000000004),
    .INIT_07(256'h000000000000101018101E000000000000000000000000000000040A11111100),
    .INIT_08(256'h0C100E0000000000000000000000000000000E1010100E000000000000000000),
    .INIT_09(256'h000000000000000000001C020C100E0000000000000000000000000000001C02),
    .INIT_0A(256'h0202020100704848487000000000000000000003020202020070484848700000),
    .INIT_0B(256'h4870000000000000000000010202020100704848487000000000000000000001),
    .INIT_0C(256'h0000000102020201007048484870000000000000000000010202020100704848),
    .INIT_0D(256'h0070083040380000000000000000000202030201004848586848000000000000),
    .INIT_0E(256'h0000000000000001010101030078406040780000000000000000000101010202),
    .INIT_0F(256'h00001E1018101E00000000000000000000000002020302010038404040380000),
    .INIT_10(256'h4078000000000000000000010202020200700830403800000000000000000000),
    .INIT_11(256'h000000000000101018101E000000000000000000000000030001020100784060),
    .INIT_12(256'h1C121C0000000000000000000000000000000E1216100C000000000000000000),
    .INIT_13(256'h000000000000000000000C121212120000000000000000000000000000001214),
    .INIT_14(256'h0303030707070707070300000000000000000000000000000000000000000000),
    .INIT_15(256'h0C0C00000000000000000000000000000C0C0C0C0C0C00000000000003030000),
    .INIT_16(256'h0F1F3B3303030F1F3B333B1F0F030300000000000C0C0C0C3C3C0C0C3C3C0C0C),
    .INIT_17(256'h3F33333F1E0C000000000000000030381C0E07030100183C3C18000000000303),
    .INIT_18(256'h0000000000000000000000000C0E070303030000000000000F1F3931333F1C1E),
    .INIT_19(256'h00000000000103070E0C0000000000000103070E0C0C0C0C0C0E070301000000),
    .INIT_1A(256'h00000000000000000003333B1F0F07070F1F3B33030000000000000C0E070301),
    .INIT_1B(256'h1C0C0C0C000000000000000000000000000000000000030303033F3F03030303),
    .INIT_1C(256'h000000000000000000000000000000000F0F0000000000000000000000003038),
    .INIT_1D(256'hC0E06070381C0E06070301000000000000000000000000000C0C000000000000),
    .INIT_1E(256'h0303030303031F0F070300000000000003070F1C3830303030381C0F07030000),
    .INIT_1F(256'h3F3F0000000000003F3F30381C0E0703000030381F0F00000000000003030303),
    .INIT_20(256'h000000003F3F30381C0E070301000000000000000F1F38300000030301000000),
    .INIT_21(256'h30381C0E07030000000000000F1F3830000000003F3F30303F3F000000000000),
    .INIT_22(256'h000000000C0C0C0C0C0E0703010000003F3F0000000000000F1F383030383F37),
    .INIT_23(256'h00000F1F383030381F0F0000000000000F1F383030381F1F303030381F0F0000),
    .INIT_24(256'h00000000000000000C0C0000000000000C0C000000000000000000000F0F0000),
    .INIT_25(256'h00000103070E1C0E0703010000000000000030381C0C0C0C000000000C0C0000),
    .INIT_26(256'h03070E1C3830000000000000000000003F3F00003F3F00000000000000000000),
    .INIT_27(256'h000000000303000003030100000030381F0F000000000030381C0E0703010001),
    .INIT_28(256'h3F3F3030303030381F0F0000000000000F1F383031333333333130381F0F0000),
    .INIT_29(256'h1F0F0000000000003F3F303030303F3F303030303F3F00000000000030303030),
    .INIT_2A(256'h3F3F303030303030303030303F3F0000000000000F1F38303030303030303038),
    .INIT_2B(256'h303030303F3F0000000000003F3F303030303F3F303030303F3F000000000000),
    .INIT_2C(256'h000000000F1F383030303030303030381F0F0000000000003030303030303F3F),
    .INIT_2D(256'h03030303030303030F0F0000000000003030303030303F3F3030303030300000),
    .INIT_2E(256'h30300000000000000F1F3930000000000000000003030000000000000F0F0303),
    .INIT_2F(256'h3F3F3030303030303030303030300000000000003030303133373E3E37333130),
    .INIT_30(256'h3E3C38303030000000000000303030303030303333373F3C3830000000000000),
    .INIT_31(256'h000000000F1F383030303030303030381F0F0000000000003030303030313337),
    .INIT_32(256'h33333030303030381F0F0000000000003030303030303F3F303030303F3F0000),
    .INIT_33(256'h1F0F0000000000003030303133373F3F303030303F3F0000000000000F1F3031),
    .INIT_34(256'h0303030303030303030303033F3F0000000000000F1F383000000F1F38303038),
    .INIT_35(256'h3830303030300000000000000F1F383030303030303030303030000000000000),
    .INIT_36(256'h000000000C1F3F3333333333303030303030000000000000030307070C0C0C18),
    .INIT_37(256'h030307070C1C18383030000000000000303038181C0F07070F1C183830300000),
    .INIT_38(256'h03030000000000003F3F30381C0E0703010000003F3F00000000000003030303),
    .INIT_39(256'h0000000000010307060E1C383060E0C000000003030303030303030303030303),
    .INIT_3A(256'h30381C0F070300000000000F0F00000000000000000000000F0F000000000000),
    .INIT_3B(256'h00003F3F00000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h303030391F0F00000000000000000000000000000000000000000003070E0C00),
    .INIT_3D(256'h00000000000000003F3F3030303030303F3F303030300000000000000F1F3930),
    .INIT_3E(256'h0F1F3830303030381F0F000000000000000000000F1F3830303030381F0F0000),
    .INIT_3F(256'h0C0C0C0E07030000000000000F1F38303F3F30381F0F00000000000000000000),
    .INIT_40(256'h070F1C1800000F1F383030381F0F000000000000000000000C0C0C0C0C0C3F3F),
    .INIT_41(256'h030303030F0F000003030000000000003030303030383C3E3733303030300000),
    .INIT_42(256'h0C0C00000F1F393000000000000000000303000000000000000000000F0F0303),
    .INIT_43(256'h0F0F030303030303030303030F0F0000000000000C0C0C0D0F0F0D0C0C0C0C0C),
    .INIT_44(256'h373300000000000000000000333333333333333F3F3C00000000000000000000),
    .INIT_45(256'h000000000F1F3830303030381F0F000000000000000000003030303030383C3E),
    .INIT_46(256'h303030381F0F000000000000303030303F3F3030303030303F3F000000000000),
    .INIT_47(256'h00000000000000003030303030383C3E3733000000000000000000000F1F3830),
    .INIT_48(256'h03070E0C0C0C0C0C0F0F0C0C0C0C0000000000003F3F00000F1F38381F0F0000),
    .INIT_49(256'h3030000000000000000000000F1F393030303030303000000000000000000000),
    .INIT_4A(256'h000000000C1F3F33333330303030000000000000000000000307070C0C1C1838),
    .INIT_4B(256'h3930303030300000000000000000000030381C0F07070F1C3830000000000000),
    .INIT_4C(256'h01000000000000003F3F1C0E070301003F3F0000000000000F1F383000000F1F),
    .INIT_4D(256'h030303030303030303030303030300000000000001030303070E1C0E07030303),
    .INIT_4E(256'h00000000000000000000000F0F01000000000000000000010F0F000000000303),
    .INIT_4F(256'h000000000000000000000018181818187E7E0000000000000000000030391F0F),
    .INIT_50(256'h3030313B1F0E000000000000000000000303000003070E1C383030381F0F0000),
    .INIT_51(256'h3F000000001818181F1F181818181F1F191D0C0E07030000000000000E1F3B31),
    .INIT_52(256'h00100B070E0C0C0E070B1000000000000000000030303030303030303030303F),
    .INIT_53(256'h0303030303030000000000000C0C0C0C0C0C3F3F000000000000000000000000),
    .INIT_54(256'h000000003F3F381C0E070303070E1C383F3F0000000003030303030303000003),
    .INIT_55(256'h3131313B1F0E000000000000000000000000000000000000000000000C0C0000),
    .INIT_56(256'h0F070000000000000303030303030363733F1E0000000000000000000E1F3B33),
    .INIT_57(256'h07070703313030303030F0F07030000000000000070F1C1830303F3F3030181C),
    .INIT_58(256'h38381C1CF8F000000000030301000000333331303030F0F07030000000000000),
    .INIT_59(256'h000000003C3C0C0C1C3830303030381F0F0000000000000007070703F1F81C1C),
    .INIT_5A(256'h0C0C06060303010100000000000000000F1F393030391F0F0303030301000000),
    .INIT_5B(256'h30000000000000000F1F38303F3F30381F0F000000000000000000003F3F1818),
    .INIT_5C(256'h00000000000000000000000303010000000000000F1F38303030303030303030),
    .INIT_5D(256'h0E000000000000000000000030303030303030303030381F0F00000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000E1F3B3131313B1F),
    .INIT_5F(256'h0000000000000000000000000C0E070300000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0E1C3933070E1C0E070301000000000000000000000000000000000000000000),
    .INIT_62(256'h03070E1C3830000000000000000000003F3F000061733F1E0000000000010307),
    .INIT_63(256'h00000000000000000000000000000000000000000C0E0733391C0E0703010001),
    .INIT_64(256'h0303030101010000010100000000000000000000000000000000000000000000),
    .INIT_65(256'h010000000000000003070E0C0C0C0C0E07030000000000000000000001030303),
    .INIT_66(256'h03070E0C3F3F0C0C3F3F0C0E07030000000000000F0F0C0E07030F0F03030303),
    .INIT_67(256'h1F0F0003070F0C0000000000030101010F010303060E0C1C1818000000000000),
    .INIT_68(256'h000000003F3F00000F1F38381F0F1C1C0F070000000000003F3F00003F3F3038),
    .INIT_69(256'h666666666773303C1F070000000000003F3F00000F1F38381F0F0003070F0C00),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000071F3C307367),
    .INIT_6B(256'h00000000001F1F0000000000000000000000000000000103070E070301000000),
    .INIT_6C(256'h6777303C1F07000000000000000000000000070F0C0C0C0F0700000000000000),
    .INIT_6D(256'h000000000000000000000000000000000F0F00000000071F3C30766666676766),
    .INIT_6E(256'h030303033F3F030303030000000000000000000000000003070E0C0E07030000),
    .INIT_6F(256'h1F1F0000000000000000000000003F3F1C0F07313F1F0000000000003F3F0000),
    .INIT_70(256'h3F3F1C0E070321303F3F0003070F0C00000000000000000000001F1F01070701),
    .INIT_71(256'h313131313F1F00003030303018181B1F1C181818181800000000000000000000),
    .INIT_72(256'h0000000000000000030707030000000000000000000000010101010101011F3F),
    .INIT_73(256'h000006060606061E0E060000000000003F3F1C0E070301003F3F0003070F0C00),
    .INIT_74(256'h0000000000000000000000000000060F1F19191F0F0600000000000000000000),
    .INIT_75(256'h0F1F3B33333333333333333B1F0F00000000000000333B1D0E070E1D3B330000),
    .INIT_76(256'h383000000C0C0000000000000F1F3B333333333B1F0F00000000000000000000),
    .INIT_77(256'h000000000F1F383030381C0E0703000003030000000000000303030303070F1C),
    .INIT_78(256'h3F3030381F0F000303010000000000003030303F3F3030381F0F0003070E0C00),
    .INIT_79(256'h190E0000000000003030303F3F3030381F0F000C0F070300000000003030303F),
    .INIT_7A(256'h3030303F3F3030381F0F00000C0C0000000000003030303F3F3030381F0F0018),
    .INIT_7B(256'h3131313B1F0F0000000000003030303F3F3030381F0F00030404030000000000),
    .INIT_7C(256'h0C0E07030F1F383030303030303030381F0F0000000000003131313131313F3F),
    .INIT_7D(256'h3E3E30303F3F000303010000000000003F3F30303E3E30303F3F0003070E0C00),
    .INIT_7E(256'h0C0C0000000000003F3F30303E3E30303F3F000C0F070300000000003F3F3030),
    .INIT_7F(256'h0F0F0303030303030F0F0003070E0C00000000003F3F30303E3E30303F3F0000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_20480x16_sub_000000_008 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_Naddra[12]_Naddr_o ),
    .dia({open_n108,open_n109,open_n110,open_n111,open_n112,open_n113,open_n114,open_n115,dia[15:8]}),
    .wea(wea),
    .doa({open_n137,open_n138,open_n139,open_n140,open_n141,open_n142,open_n143,open_n144,inst_doa_i0_015,inst_doa_i0_014,inst_doa_i0_013,inst_doa_i0_012,inst_doa_i0_011,inst_doa_i0_010,inst_doa_i0_009,inst_doa_i0_008}));
  // address_offset=4096;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=16;working_depth=4096;working_width=8;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'hC0C000C0C080000000000000C0C0000000000000C0C0000080C0C00000000000),
    .INIT_01(256'h00000000C0C0000000000000C0C00000C0C0000000000000C0C0000000000000),
    .INIT_02(256'hB030303030300000C060600000000000C0E070303030303030303070E0C00000),
    .INIT_03(256'h80C0C00000000000C0F0303030303030F0C0000000000000000000003070F0F0),
    .INIT_04(256'hC0F0303030303030F0C000C0C080000000000000C0F0303030303030F0C00000),
    .INIT_05(256'hF0C00000C0C0000000000000C0F0303030303030F0C00000C060600000000000),
    .INIT_06(256'h000000002070E0C08080C0E0702000000000000000000000C0F0303030303030),
    .INIT_07(256'h30303030303000000000000000000000C0E070303030303030B0B070E0D00000),
    .INIT_08(256'hC080000000000000C0E07030303030303030000080C0C00000000000C0E07030),
    .INIT_09(256'hC0E070303030303030300000C0C0000000000000C0E0703030303030303000C0),
    .INIT_0A(256'h70E0C0000000000000000000000000000080C0E07030000080C0C00000000000),
    .INIT_0B(256'h000000000080C0C0C0C08000008080800000000000000000000000C0E0703030),
    .INIT_0C(256'h7070F0F0B030000080C0C0000000000030B0F0F07070F0F0B030000000000000),
    .INIT_0D(256'hC06060000000000030B0F0F07070F0F0B03000C0C08000000000000030B0F0F0),
    .INIT_0E(256'h30B0F0F07070F0F0B0300000C0C000000000000030B0F0F07070F0F0B0300000),
    .INIT_0F(256'hF8F00000000000000000000030B0F0F07070F0F0B03000008080000000000000),
    .INIT_10(256'h00000000C0C0000000000000C0C000000000000000000000F8F88080FCFC8C9C),
    .INIT_11(256'hF0F03070E0C0000080C0C00000000000E0E00000F0F03070E0C0000000000000),
    .INIT_12(256'hC0C0000000000000E0E00000F0F03070E0C000C0C080000000000000E0E00000),
    .INIT_13(256'hC0C0000000000000000000000000000000000000E0E00000F0F03070E0C00000),
    .INIT_14(256'h000000C0C080000000000000C0C00000000000000000000080C0C00000000000),
    .INIT_15(256'h00000000C0C000000000000000000000C0C0000000000000C0C0000000000000),
    .INIT_16(256'h30303070E0C00000C060600000000000C0E070303030F0E06060C0F080800000),
    .INIT_17(256'h80C0C00000000000C0E0703030303070E0C00000000000000000000030303030),
    .INIT_18(256'hC0E0703030303070E0C000C0C080000000000000C0E0703030303070E0C00000),
    .INIT_19(256'hE0C00000C0C0000000000000C0E0703030303070E0C00000C060600000000000),
    .INIT_1A(256'h00000000000000000000F0F0000000000000000000000000C0E0703030303070),
    .INIT_1B(256'h70303030303000000000000000000000C0E070303030B070E0D0000000000000),
    .INIT_1C(256'hC08000000000000030B0F0F0703030303030000080C0C0000000000030B0F0F0),
    .INIT_1D(256'h30B0F0F07030303030300000C0C000000000000030B0F0F070303030303000C0),
    .INIT_1E(256'hC080000000000000C0E07030303030B0F0F070303030000080C0C00000000000),
    .INIT_1F(256'hC0E07030303030B0F0F0703030300000C0C00000000000000000000080C0C0C0),
    .INIT_20(256'h8686868E9C98FEFEFCF880800000F8F818189898989898989898FEFEFCF88080),
    .INIT_21(256'hE0C0000000006060606060E0C080F8FC8E86C0E0E0C000000000F8F8181C8E86),
    .INIT_22(256'h1C3870E0C080F8FC8E86C0E0E0C000000000060E1C3870E0C080FEFE8080C0E0),
    .INIT_23(256'hE0E0E0C08000000000006060606060E0C68EFCF88080C0E0E0C000000000060E),
    .INIT_24(256'h00008080C0C0E0E0F0FCFEFCF0E0E0C0C0808000000000C08098BCFEFEFEFCD8),
    .INIT_25(256'hFEFEFCF8F0E0E0C08080000000000080C0C0E0F0F8FCFEFEFE7E3C1800000000),
    .INIT_26(256'h00000000000000000000C0E070303070E0C0000000000000000000C08098BCFE),
    .INIT_27(256'hE0F8381C0C0C0C0C1C38F8E000000000000000000000C0E0F0F0F0F0E0C00000),
    .INIT_28(256'h808080000000000000000000E0F8F8FCFCFCFCFCFCF8F8E00000000000000000),
    .INIT_29(256'h00000080C0E0F0F0F8F8F0F0E0C0800000000000000000001030E0E0C0E0F8FC),
    .INIT_2A(256'hFEFEFE9E9E9EFCFCF8E000000000E0F8FC3CCEF6FEFEFE9E9E9EFCFCF8E00000),
    .INIT_2B(256'hF8E000000000E0F8FCFCFEF6CE3EFE9E9E9EFCFCF8E000000000E0F8FCFCFE06),
    .INIT_2C(256'hFC3CCE763E3E7E9E9E9EFCFCF8E000000000E0F8FC3CCEF6FEFEFEFE8EFEFCFC),
    .INIT_2D(256'h8EFEFCFCF8E000000000E0F83CDC5EDE0EF6FE9E9E9EFCFCF8E000000000E0F8),
    .INIT_2E(256'h0000E01804C4320A020202626262040418E000000000E0F83CDC5EDE0EF6FEFE),
    .INIT_2F(256'h32C202626262040418E000000000E018040402FA020202626262040418E00000),
    .INIT_30(256'h18E000000000E01804C4320A020202027202040418E000000000E0180404020A),
    .INIT_31(256'hC424A222F20A02626262040418E000000000E01804C4328AC2C2826262620404),
    .INIT_32(256'h1404FC00000000000000E018C424A222F20A02027202040418E000000000E018),
    .INIT_33(256'h000000000000C020900804089020C00000000000000000000000FC0414A444A4),
    .INIT_34(256'h86E6E6868E1C38F0E00000000000000040407048700000000000000000000000),
    .INIT_35(256'hE0000000000000E0F0381C0E060606060E1C38F0E0000000000000E0F0381C8E),
    .INIT_36(256'h3C7E666666666666666666667E3C0000000000E0F0381CCEE6E6E6E6CE1C38F0),
    .INIT_37(256'h666666667E3C0000000000000C0C0C0C0C0C0C0C0C0C7C3C1C0C000000000000),
    .INIT_38(256'h000000000C0C0C0C0C0C0C0C0C0C7C3C1C0C0000000000003C7E666666666666),
    .INIT_39(256'h0C0C0C0C0C0C7C3C1C0C0000000000003C7E666666666666666666667E3C0000),
    .INIT_3A(256'h000000000000000000000000000000000000000000000000000000000C0C0C0C),
    .INIT_3B(256'h3C7E666666666666666666667E3C000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000C0C0C0C0C0C0C0C0C0C7C3C1C0C000000000000),
    .INIT_3D(256'h0000000042422418182442420000000000000000000000004242241818244242),
    .INIT_3E(256'h0000808080808080808000000000000000000000000080C0E06060E0C0800000),
    .INIT_3F(256'hF0E0000000000000000000000000F0F000C0E070F0E000000000000000000000),
    .INIT_40(256'h000000000000C0C0F0F0C0C0C0C0000000000000000000000000E0F070E0E070),
    .INIT_41(256'h30F0E000E0E0000000000000000000000000E0F030F0E000F0F0000000000000),
    .INIT_42(256'h00000000000000000000808080C0E070F0F0000000000000000000000000E0F0),
    .INIT_43(256'h0000E0F030F0F030F0E0000000000000000000000000E0F030F0E030F0E00000),
    .INIT_44(256'hFE0000000000000000F0F00000F0F00000F0F000000000000000000000000000),
    .INIT_45(256'hFE06060606F6F606060606FEFE000000000000FEFE06868686F6F686868606FE),
    .INIT_46(256'h060606FEFE000000000000FEFE060686C6E070381C0E06E0E0000000000000FE),
    .INIT_47(256'h000000FEFE063676E6C6C6E6763606FEFE000000000000FEFE06060606060606),
    .INIT_48(256'hF0F03070E0C0000000000000000000FCFC0C8C8CCCCC0CFCFC181838F0E08000),
    .INIT_49(256'h0000000000000000C0E07070E0E07070E0C00000000000000000000030303030),
    .INIT_4A(256'hC0E0703030303070E0C000000000000000000000C0E0703000003070E0C00000),
    .INIT_4B(256'hF0F000000000000000000000F0F00000C0C00000F0F000000000000000000000),
    .INIT_4C(256'h00000000E0F03030F0F00000C0C00000000000000000000000000000C0C00000),
    .INIT_4D(256'h00000000C0C00000000000000000000030303030F0F030303030000000000000),
    .INIT_4E(256'h00000000000000000080C0C0C0C0C0C0F0F000000000000000000000C0C00000),
    .INIT_4F(256'hF0F00000000000000000000000000000000000003070E0C08080C0E070300000),
    .INIT_50(256'h3030000000000000000000003030303030B0F0F0703000000000000000000000),
    .INIT_51(256'h00000000C0E0703030303070E0C0000000000000000000003070F0F0B0303030),
    .INIT_52(256'hB0303070E0C00000000000000000000000000000C0E07070E0C0000000000000),
    .INIT_53(256'h0000000000000000C0C08000C0E07070E0C0000000000000000000003070E0C0),
    .INIT_54(256'h0000000000000000F0F000000000000000000000C0E07030F0F00000F0F00000),
    .INIT_55(256'h303000000000000000000000C0E0703030303030303000000000000000000000),
    .INIT_56(256'h00000000C0E07030303030303030000000000000000000000080C0E070303030),
    .INIT_57(256'h0080C0E07030000000000000000000003070E0C08080C0E07030000000000000),
    .INIT_58(256'h3030000000000000F0F000000080C0E0F0F00000000000000000000000000000),
    .INIT_59(256'hF0F030303030F0F030303030F0F000000000000000008080C0C0C0E0E0607030),
    .INIT_5A(256'h0000000000000000000000006060C0C080800000000000000000000000000000),
    .INIT_5B(256'h00000018BCBC180000000080C0E06000000000000000000000008080C0C06060),
    .INIT_5C(256'h0000B0F0703070F0B00000000000000078404040400000000000000000000000),
    .INIT_5D(256'hE0E0000000000000000000000000E0F03030F0E0000000000000000000000000),
    .INIT_5E(256'h000000000000F0F03030F0F03030000000000000000000000000E0E000000000),
    .INIT_5F(256'h00C00030F0E0000000000000000000000000E0E000E0F030F0E0000000000000),
    .INIT_60(256'h000000000000000000E0F03030F0F030F0E00000000000000000000000000000),
    .INIT_61(256'h00008080808080008080000000000000000000000000303030F0E00000000000),
    .INIT_62(256'hC0000000000000000000000000C0E06060E0E000606000000000000000000000),
    .INIT_63(256'h000000000000C0C00000000000000000000000000000000000003070E0C080C0),
    .INIT_64(256'h3030F0E0000000000000000000000000000018989898F8F00000000000000000),
    .INIT_65(256'h00000000000000000000C0E0703070E0C0000000000000000000000000003030),
    .INIT_66(256'h003030F0F03030F0F00000000000000000000000000000E0F03030F0E0000000),
    .INIT_67(256'hE0C00000000000000000000000000000000060E0C00000000000000000000000),
    .INIT_68(256'h000000000000C0C00000C0C00000000000000000000000000000C0E060E0C000),
    .INIT_69(256'hE07030303000000000000000000000000000E0F0303030303000000000000000),
    .INIT_6A(256'h0000000000000000000060F0B8989818180000000000000000000000000080C0),
    .INIT_6B(256'h00C0E06060E0E06060600000000000000000000000003070E0C0E07030000000),
    .INIT_6C(256'h0000000000000000000000000000E0E00080C0E0E0E000000000000000000000),
    .INIT_6D(256'h00F8F8787818187878F8F800000000000000000000E0F0B818383818B8F0E000),
    .INIT_6E(256'h78F0E000000000000000000000F8F8F8F81818F8F8F8F8000000000000000000),
    .INIT_6F(256'h0000000000E0F0F8F81818F8F8F0E000000000000000000000E0F07878181878),
    .INIT_70(256'h0080808080808080808080800000000000000000008080000000000000000000),
    .INIT_71(256'h80808080000000000000000000FFFF0000000000000000000000000000000000),
    .INIT_72(256'h80808080808080000000000000000000000000000000000000FFFF8080808080),
    .INIT_73(256'h0000000000000000808080808080808080808080808080808080808080808080),
    .INIT_74(256'h808080808080808080FFFF808080808080808080808080808080808080FFFF00),
    .INIT_75(256'h0080808080808080808080800000000000000000008080000000000000000000),
    .INIT_76(256'h80808080000000000000000000FFFF0000000000000000000000000000000000),
    .INIT_77(256'h80808080808080000000000000000000000000000000000000FFFF8080808080),
    .INIT_78(256'h0000000000000000808080808080808080808080808080808080808080808080),
    .INIT_79(256'h808080808080808080FFFF808080808080808080808080808080808080FFFF00),
    .INIT_7A(256'hC040404040404040404040400000000000000000C04040C00000000000000000),
    .INIT_7B(256'h404040400000000000000000FF0000FF00000000000000000000000000000000),
    .INIT_7C(256'h404040404040404000000000000000000000000000000000FF00007F40404040),
    .INIT_7D(256'h0000000000000000404040404040404040404040404040404040404040404040),
    .INIT_7E(256'h40404040404040407F00007F404040404040404040404040404040407F0000FF),
    .INIT_7F(256'hC040404040404040404040400000000000000000C04040C00000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_20480x16_sub_004096_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_addra[12]_Naddra_o ),
    .dia({open_n165,open_n166,open_n167,open_n168,open_n169,open_n170,open_n171,open_n172,dia[7:0]}),
    .wea(wea),
    .doa({open_n194,open_n195,open_n196,open_n197,open_n198,open_n199,open_n200,open_n201,inst_doa_i1_007,inst_doa_i1_006,inst_doa_i1_005,inst_doa_i1_004,inst_doa_i1_003,inst_doa_i1_002,inst_doa_i1_001,inst_doa_i1_000}));
  // address_offset=4096;data_offset=8;depth=4096;width=8;num_section=1;width_per_section=8;section_size=16;working_depth=4096;working_width=8;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0F0F000C0F070300000000000F0F0303030303030F0F00030301000000000000),
    .INIT_01(256'h000000000F0F0303030303030F0F00000C0C0000000000000F0F030303030303),
    .INIT_02(256'h33373E3C38300018190E0000000000003F3F303030307C7C303030303F3F0000),
    .INIT_03(256'h03010000000000000F3F3030303030303F0F0003070E0C000000000030303031),
    .INIT_04(256'h0F3F3030303030303F0F000C0F070300000000000F3F3030303030303F0F0003),
    .INIT_05(256'h3F0F00000C0C0000000000000F3F3030303030303F0F0018190E000000000000),
    .INIT_06(256'h0000000010381C0F07070F1C3810000000000000000000000F3F303030303030),
    .INIT_07(256'h3030303030300003070E0C00000000002F1F383434323231313030381F0F0000),
    .INIT_08(256'h0F070300000000000F1F3830303030303030000303010000000000000F1F3830),
    .INIT_09(256'h0F1F383030303030303000000C0C0000000000000F1F3830303030303030000C),
    .INIT_0A(256'h0C0F0F0C3F3F0000000000000303030303070F1C383000030301000000000000),
    .INIT_0B(256'h003030303737313030313737333B191D0F060000000000003F3F0C0F0F0C0C0C),
    .INIT_0C(256'h303030391F0F000303010000000000000F1F3930303030391F0F0003070E0C00),
    .INIT_0D(256'h190E0000000000000F1F3930303030391F0F000C0F070300000000000F1F3930),
    .INIT_0E(256'h0F1F3930303030391F0F00000C0C0000000000000F1F3930303030391F0F0018),
    .INIT_0F(256'h1F1F000000000000000000000F1F3930303030391F0F00030404030000000000),
    .INIT_10(256'h0C0E07030F1F3830303030381F0F000000000000000000000F1F39391F0F0101),
    .INIT_11(256'h3F3F30381F0F000303010000000000000F1F38303F3F30381F0F0003070E0C00),
    .INIT_12(256'h0C0C0000000000000F1F38303F3F30381F0F000C0F070300000000000F1F3830),
    .INIT_13(256'h0F0F0303030303030F0F0003070E0C00000000000F1F38303F3F30381F0F0000),
    .INIT_14(256'h0F0F000C0F070300000000000F0F0303030303030F0F00030301000000000000),
    .INIT_15(256'h000000000F0F0303030303030F0F00000C0C0000000000000F0F030303030303),
    .INIT_16(256'h30383C3E37330018190E0000000000000F1F383030381F0F0000030001010000),
    .INIT_17(256'h03010000000000000F1F3830303030381F0F0003070E0C000000000030303030),
    .INIT_18(256'h0F1F3830303030381F0F000C0F070300000000000F1F3830303030381F0F0003),
    .INIT_19(256'h1F0F00000C0C0000000000000F1F3830303030381F0F0018190E000000000000),
    .INIT_1A(256'h000000000000030300003F3F0000030300000000000000000F1F383030303038),
    .INIT_1B(256'h3030303030300003070E0C00000000002F1F3834323130381F0F000000000000),
    .INIT_1C(256'h0F070300000000000F1F3930303030303030000303010000000000000F1F3930),
    .INIT_1D(256'h0F1F393030303030303000000C0C0000000000000F1F3930303030303030000C),
    .INIT_1E(256'h313F3F30303030000F1F383000000F1F39303030303000030301000000000000),
    .INIT_1F(256'h0F1F383000000F1F39303030303000000C0C0000000000303030303F3F313030),
    .INIT_20(256'h6161617139197F7F3F1F010100001F1F181819191919191919197F7F3F1F0101),
    .INIT_21(256'h07030000000006060606060703011F3F716103070703000000001F1F18387161),
    .INIT_22(256'h0606060763713F1F010103070703000000006070381C0E0703017F7F01010307),
    .INIT_23(256'h070707030100000000006070381C0E0703011F3F716103070703000000000606),
    .INIT_24(256'h00000101030307070F3F7F3F0F070703030101000000000301193D7F7F7F3F1B),
    .INIT_25(256'h7F7F3F1F0F07070301010000000000010303070F1F3F7F7F7F7E3C1800000000),
    .INIT_26(256'h0000000000000000000003070E0C0C0E07030000000000000000000301193D7F),
    .INIT_27(256'h071F1C3830303030381C1F070000000000000000000003070F0F0F0F07030000),
    .INIT_28(256'h030303010100000000000000071F1F3F3F3F3F3F3F1F1F070000000000000000),
    .INIT_29(256'h00001C0703010000000000000103071C000000000000000010180E0F070F3F7F),
    .INIT_2A(256'h7F7F7F7979793F3F1F0700000000071F3F3C736F7F7F7F7979793F3F1F070000),
    .INIT_2B(256'h1F0700000000071F3F3F7F6F737C7F7979793F3F1F0700000000071F3F3F7F60),
    .INIT_2C(256'h3F3C736E7C7C7E7979793F3F1F0700000000071F3F3C736F7F7F7F7979793F3F),
    .INIT_2D(256'h79793F3F1F0700000000071F3C3B7B7A706F7F7979793F3F1F0700000000071F),
    .INIT_2E(256'h0000071820234C504040404646462020180700000000071F3C3B7B7A706F7F79),
    .INIT_2F(256'h4C4340464646202018070000000007182020405F404040464646202018070000),
    .INIT_30(256'h180700000000071820234C504040404646462020180700000000071820204050),
    .INIT_31(256'h232444454F50404646462020180700000000071820234C514343414646462020),
    .INIT_32(256'h090403000000000000000718232444454F504046464620201807000000000718),
    .INIT_33(256'h0000000000003F202825222528203F0000000000000000000000030409102010),
    .INIT_34(256'h6167676171381C0F07000000000000000000000000000E010608070000000000),
    .INIT_35(256'h07000000000000070F1C38706060606070381C0F07000000000000070F1C3871),
    .INIT_36(256'h3C7E666666666666666666667E3C0000000000070F1C38736767676773381C0F),
    .INIT_37(256'h0C0C7C3C1C0C0000000000003C7E666666666666666666667E3C000000000000),
    .INIT_38(256'h000000000C0C0C0C0C0C0C0C0C0C7C3C1C0C0000000000000C0C0C0C0C0C0C0C),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h1C0C0000000000003C7E666666666666666666667E3C00000000000000000000),
    .INIT_3B(256'h42422418182442420000000000000000000000000C0C0C0C0C0C0C0C0C0C7C3C),
    .INIT_3C(256'h666666667E3C0000000000004242241818244242000000000000000000000000),
    .INIT_3D(256'h000000000C0C0C0C0C0C0C0C0C0C7C3C1C0C0000000000003C7E666666666666),
    .INIT_3E(256'h0000010101010107030100000000000000000000000001030706060703010000),
    .INIT_3F(256'h07070000000000000000000000000F0F0703010C0F0700000000000000000000),
    .INIT_40(256'h00000000000000000F0F06030100000000000000000000000000070700010100),
    .INIT_41(256'h0C0F0F0E0703000000000000000000000000070F000F0F0C0F0F000000000000),
    .INIT_42(256'h000000000000000000000101010100000F0F000000000000000000000000070F),
    .INIT_43(256'h0000070700070F0C0F07000000000000000000000000070F0C0F070C0F070000),
    .INIT_44(256'h7F00000000000000000F0F00000F0F00000F0F00000000000000000000000000),
    .INIT_45(256'h7F606060606F6F606060607F7F0000000000007F7F606161616F6F616161607F),
    .INIT_46(256'h6060607F7F0000000000007F7F60606163676E6C6060607F7F0000000000007F),
    .INIT_47(256'h0000007F7F606C6E676363676E6C607F7F0000000000007F7F60606060606060),
    .INIT_48(256'h3F3F30381F0F0000000000000000003F3F3031313333303F3F18181C0F070100),
    .INIT_49(256'h00000000000000003F3F30303F3F30303F3F0000000000000000000030303030),
    .INIT_4A(256'h3F3F3030303030303F3F000000000000000000000F1F3830303030381F0F0000),
    .INIT_4B(256'h3F3F000000000000000000003F3F30303F3F30303F3F00000000000000000000),
    .INIT_4C(256'h000000000F1F3830303030381F0F00000000000000000000303030303F3F3030),
    .INIT_4D(256'h030303030F0F00000000000000000000303030303F3F30303030000000000000),
    .INIT_4E(256'h00000000000000000F1F3930000000000303000000000000000000000F0F0303),
    .INIT_4F(256'h3F3F303030303030303000000000000000000000303030313F3F313030300000),
    .INIT_50(256'h3830000000000000000000003030303033373F3C383000000000000000000000),
    .INIT_51(256'h000000000F1F3830303030381F0F000000000000000000003030303133373E3C),
    .INIT_52(256'h333330381F0F00000000000000000000303030303F3F30303F3F000000000000),
    .INIT_53(256'h0000000000000000303133373F3F30303F3F000000000000000000000F1F3831),
    .INIT_54(256'h03030303030303033F3F000000000000000000003F3F00003F3F30381F0F0000),
    .INIT_55(256'h3030000000000000000000000F1F383030303030303000000000000000000000),
    .INIT_56(256'h000000003F3F33333333303030300000000000000000000003070F1C38303030),
    .INIT_57(256'h03070F1C38300000000000000000000030381C0F07070F1C3830000000000000),
    .INIT_58(256'h30300000000000003F3F1C0E070301003F3F0000000000000000000003030303),
    .INIT_59(256'h3F3F000000003F3F000000003F3F000000000000030307070C0C0C1F1F183830),
    .INIT_5A(256'h00000000000000000000000018180C0C07070303000000000000000000000000),
    .INIT_5B(256'h00000003076773381C0E0703317878300000000000000000030307070C0C1818),
    .INIT_5C(256'h0000070F0C0C0C0F070000000000000000000000000009090B0D090000000000),
    .INIT_5D(256'h0F070000000000000000000000000F0F0C0C0F0F0C0C00000000000000000000),
    .INIT_5E(256'h000000000000070F0C0C0F070000000000000000000000000000070F0C0C0C0C),
    .INIT_5F(256'h030F03030301000000000000000000000000070F0C0F0F0C0F07000000000000),
    .INIT_60(256'h000000000000000000070F0C00070F0C0F070000000000000000000000000303),
    .INIT_61(256'h000001010103030001010000000000000000000000000C0C0C0F0F0C0C0C0000),
    .INIT_62(256'h0C0C000000000000000000000003070600000000000000000000000000000000),
    .INIT_63(256'h00000000000001030303030303030000000000000000000000000C0C0C0F0F0D),
    .INIT_64(256'h0C0C0F0F0000000000000000000000000000181919191F1F0000000000000000),
    .INIT_65(256'h0000000000000000000003070E0C0E0703000000000000000000000000000C0C),
    .INIT_66(256'h000000070F0C0C0F070000000000000000000000000C0C0F0F0C0C0F0F000000),
    .INIT_67(256'h0F070000000000000000000000000C0C0C0C0E0F0D0000000000000000000000),
    .INIT_68(256'h000000000000010303030F0F0303000000000000000000000000070F00070F0C),
    .INIT_69(256'h070E0C0C0C00000000000000000000000000070F0C0C0C0C0C00000000000000),
    .INIT_6A(256'h00000000000000000000060F1D19191818000000000000000000000000000103),
    .INIT_6B(256'h000307060001030706060000000000000000000000000C0E0703070E0C000000),
    .INIT_6C(256'h00000000000000000000000000000F0F070301000F0F00000000000000000000),
    .INIT_6D(256'h001F1F1E1E18181E1E1F1F00000000000000000000070F1D181C1C181D0F0700),
    .INIT_6E(256'h1E0F07000000000000000000001F1F1F1F18181F1F1F1F000000000000000000),
    .INIT_6F(256'h0000000000070F1F1F18181F1F0F0700000000000000000000070F1E1E18181E),
    .INIT_70(256'h0001010101010101010101010000000000000000000101000000000000000000),
    .INIT_71(256'h0101010100000000000000000001010000000000000000000000000000000000),
    .INIT_72(256'h0101010101010100000000000000000000000000000000000001010101010101),
    .INIT_73(256'h0000000000000000010101010101010101010101010101010101010101010101),
    .INIT_74(256'h0101010101010101010101010101010101010101010101010101010101010100),
    .INIT_75(256'h00FFFF010101010101010101000000000000000000FFFF000000000000000000),
    .INIT_76(256'h01010101000000000000000000FFFF0000000000000000000000000000000000),
    .INIT_77(256'h0101010101FFFF000000000000000000000000000000000000FFFF0101010101),
    .INIT_78(256'h0000000000000000010101010101010101FFFF01010101010101010101010101),
    .INIT_79(256'h010101010101010101FFFF010101010101010101010101010101010101FFFF00),
    .INIT_7A(256'h0302020202020202020202020000000000000000030202030000000000000000),
    .INIT_7B(256'h0202020200000000000000000302020300000000000000000000000000000000),
    .INIT_7C(256'h0202020202020202000000000000000000000000000000000302020202020202),
    .INIT_7D(256'h0000000000000000020202020202020202020202020202020202020202020202),
    .INIT_7E(256'h0202020202020202020202020202020202020202020202020202020202020203),
    .INIT_7F(256'hFF0000FE02020202020202020000000000000000FF0000FF0000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_20480x16_sub_004096_008 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_addra[12]_Naddra_o ),
    .dia({open_n222,open_n223,open_n224,open_n225,open_n226,open_n227,open_n228,open_n229,dia[15:8]}),
    .wea(wea),
    .doa({open_n251,open_n252,open_n253,open_n254,open_n255,open_n256,open_n257,open_n258,inst_doa_i1_015,inst_doa_i1_014,inst_doa_i1_013,inst_doa_i1_012,inst_doa_i1_011,inst_doa_i1_010,inst_doa_i1_009,inst_doa_i1_008}));
  // address_offset=8192;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=16;working_depth=4096;working_width=8;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h404040400000000000000000FF0000FF00000000000000000000000000000000),
    .INIT_01(256'h40404040404040C000000000000000000000000000000000FF00007F40404040),
    .INIT_02(256'h0000000000000000404040404040404040404040404040404040404040404040),
    .INIT_03(256'h40404040404040407F00007F404040404040404040404040404040407F0000FF),
    .INIT_04(256'hC0C0C0C0C0C0C0C0C0C0C0C00000000000000000C0C0C0C00000000000000000),
    .INIT_05(256'hC0C0C0C00000000000000000FFFFFFFF00000000000000000000000000000000),
    .INIT_06(256'hC0C0C0C0C0C0C0C000000000000000000000000000000000FFFFFFFFC0C0C0C0),
    .INIT_07(256'h0000000000000000C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0),
    .INIT_08(256'hC0C0C0C0C0C0C0C0FFFFFFFFC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0FFFFFFFF),
    .INIT_09(256'hC0C0C0C0C0C0C0C0C0C0C0C00000000000000000C0C0C0C00000000000000000),
    .INIT_0A(256'hC0C0C0C00000000000000000FFFFFFFF00000000000000000000000000000000),
    .INIT_0B(256'hC0C0C0C0C0C0C0C000000000000000000000000000000000FFFFFFFFC0C0C0C0),
    .INIT_0C(256'h0000000000000000C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0),
    .INIT_0D(256'hC0C0C0C0C0C0C0C0FFFFFFFFC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0FFFFFFFF),
    .INIT_0E(256'h8000008080808000008080804040400000404040400000404040400000404040),
    .INIT_0F(256'h00000000C0C0C00000C0C0C0C00000C0C0C0C00000C0C0C08080800000808080),
    .INIT_10(256'h0000000000737300000000000000000000000000000000007300007300000000),
    .INIT_11(256'h4040404040404040000000000000000073737373000000000000000000000000),
    .INIT_12(256'h40404040404040404040404040404040404040404040404040404040407F7F40),
    .INIT_13(256'hFF0000FF00000000000000000000000000000000FF0000FF8080808080808080),
    .INIT_14(256'hC0C0C0C0C0C0C0C0C0C0C0C0FFFFFFFF80808080808080808080808080808080),
    .INIT_15(256'h80808080FFFFFFFFC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0FFFFFFFFC0C0C0C0),
    .INIT_16(256'h8080808080808080C0C0C0C0C0C0C0C0C0FFFFC0C0C0C0C0C0C0C0C080808080),
    .INIT_17(256'hC0C0C0C0C0C0C0C0C0FFFFC0C0C0C0C0C0C0C0C08080808080808080FFFFFFFF),
    .INIT_18(256'hFFFFFFFF8080808080808080000000000000000000FFFFC0C0C0C0C0C0C0C0C0),
    .INIT_19(256'h00000000C0C0C0C0C0C0C0C0C0FFFF0000000000000000000000000000000000),
    .INIT_1A(256'h0000000000C0C0C0C0C0C0C0C0C0C0C08080808080808080FFFFFFFF00000000),
    .INIT_1B(256'h0000000000000000000000000000000080808080808080808080808000000000),
    .INIT_1C(256'h8080808080808080808080800000000000000000C0C0C0C0C0C0C0C0C0C0C000),
    .INIT_1D(256'hFFFFFFFF8080808080808080C0C0C0C0C0C0C0C0C0FFFFC0C0C0C0C0C0C0C0C0),
    .INIT_1E(256'h80808080C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C08080808080808080),
    .INIT_1F(256'h00000000FFFFFFFF808080808080808080808080808080808080808080808080),
    .INIT_20(256'h0000000000000000000000000000000000FFFFC0C0C0C0C0C0C0C0C000000000),
    .INIT_21(256'hC0C0C0C0C0C0C0C0C0FFFF0000000000000000008080808080808080FFFFFFFF),
    .INIT_22(256'hFFFFFFFF40404040404040400000000000000000FFC0C0FFC0C0C0C0C0C0C0C0),
    .INIT_23(256'h00000000C0C0C0C0C0C0C0C0FFC0C0FF00000000000000000000000000000000),
    .INIT_24(256'h00000000C0C0C0C0C0C0C0C0C0C0C0C04040404040404040FFFFFFFF00000000),
    .INIT_25(256'h00000000000000000000000000000000C0C0C0C0404040404040404000000000),
    .INIT_26(256'h4040404040404040C0C0C0C00000000000000000C0C0C0C0C0C0C0C0C0C0C0C0),
    .INIT_27(256'h7F7F7F7F4040404040404040C0C0C0C0C0C0C0C0FFC0C0FFC0C0C0C0C0C0C0C0),
    .INIT_28(256'h404040404040404040404040FFFFFFFFC0C0C0C0C0C0C0C04040404040404040),
    .INIT_29(256'hC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0FFFFFFFF40404040),
    .INIT_2A(256'hC0C0C0C0C0C0C0C04040404040404040404040404040404040404040C0C0C0C0),
    .INIT_2B(256'hC0C0C0C0C0C0C0C0C0C0C0C040404040404040404040404040404040C0C0C0C0),
    .INIT_2C(256'hFFC0C0FFC0C0C0C0C0C0C0C04040404040404040FFFFFFFFC0C0C0C0C0C0C0C0),
    .INIT_2D(256'hC0C0C0C0C0C0C0C0C0C0C0C0FFFFFFFF40404040404040404040404040404040),
    .INIT_2E(256'h40404040FFFFFFFFC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0FFFFFFFFC0C0C0C0),
    .INIT_2F(256'hC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0FFC0C0FFC0C0C0C0C0C0C0C040404040),
    .INIT_30(256'h40404040404040407F7F7F7F4040404040404040C0C0C0C0C0C0C0C0FF0000FF),
    .INIT_31(256'hFFFFFFFF40404040404040400000000000000000FF0000FFC0C0C0C0C0C0C0C0),
    .INIT_32(256'hC0C0C0C00000000000000000FFC0C0FFC0C0C0C0C0C0C0C00000000000000000),
    .INIT_33(256'hC0C0C0C0FFFFFFFF00000000000000000000000000000000FFFFFFFFC0C0C0C0),
    .INIT_34(256'h0000000000000000C0C0C0C0C0C0C0C0FFC0C0FF0000000000000000C0C0C0C0),
    .INIT_35(256'hC0C0C0C0C0C0C0C0FF0000FF00000000000000004040404040404040FFFFFFFF),
    .INIT_36(256'hFFFFFFFF4040404040404040C0C0C0C0C0C0C0C0FFC0C0FF4040404040404040),
    .INIT_37(256'h000000000000000000000000FF0000FF0000000000000000C0C0C0C0C0C0C0C0),
    .INIT_38(256'hC0C0C0C0C0C0404040404040404040400000000000000000FFFFFFFF00000000),
    .INIT_39(256'h808080808080808040404040404040404040C0C0C0C0C0C0C0C0C0C0C0C0C0C0),
    .INIT_3A(256'h80808080808080808080808080808080808080808080808080808080FF8080FF),
    .INIT_3B(256'h40FFFF000000000000000000000000000000000000FFFF404040404040404040),
    .INIT_3C(256'hFFFFFFFF7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F4040404040404040),
    .INIT_3D(256'h7F7F7F7F7F00007F7F7F7F7F7F7F7F7FFFFFFFFFFFFFFFFFFF0000FFFFFFFFFF),
    .INIT_3E(256'h40404040404040407F7F7F7F7F7F7F7F7F0000FF00000000000000007F7F7F7F),
    .INIT_3F(256'h0000000000000000FF00007F7F7F7F7F7F7F7F7F404040404040404040404040),
    .INIT_40(256'h7F00007F404040404040404040404040404040407F00007F7F7F7F7F7F7F7F7F),
    .INIT_41(256'h000000007F7F7F7F7F7F7F7F7F0000FF00000000000000007F7F7F7F7F7F7F7F),
    .INIT_42(256'h4040404040404040404040404040404040404040404040407F0000FF00000000),
    .INIT_43(256'h4040404040404040404040404040404040404040404040404040404040404040),
    .INIT_44(256'h0000000000000000FF00007F7F7F7F7F7F7F7F7F0000000000000000FF00007F),
    .INIT_45(256'h7F00007F404040404040404040404040404040407F00007F7F7F7F7F7F7F7F7F),
    .INIT_46(256'hFFFFFFFF7F7F7F7F7F7F7F7F7F0000FFFFFFFFFFFFFFFFFF7F7F7F7F7F7F7F7F),
    .INIT_47(256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F40404040404040407F0000FFFFFFFFFF),
    .INIT_48(256'h40404040404040407F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F),
    .INIT_49(256'hFFFFFFFFFFFFFFFFFF00007F7F7F7F7F7F7F7F7FFFFFFFFFFFFFFFFFFF00007F),
    .INIT_4A(256'hFF00007F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F0000FF0000000000000000),
    .INIT_4B(256'h000000000000000000000000C040404040404040404040400000000000000000),
    .INIT_4C(256'h404040407F0000FFFFFFFFFFFFFFFFFF4040404040404040404040C000000000),
    .INIT_4D(256'h7F7F7F7F7F7F7F7FFFFFFFFFFFFFFFFFFF00007F404040404040404040404040),
    .INIT_4E(256'h7F7F7F7F7F7F7F7F7F7F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F),
    .INIT_4F(256'hFF00007F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F0000FFFFFFFFFFFFFFFFFF),
    .INIT_50(256'hFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F7F7F7F7F7F7F7F7FFFFFFFFFFFFFFFFF),
    .INIT_51(256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7FFFFFFFFFFF),
    .INIT_52(256'h000000000000000040404040404040404040404040404040404040407F7F7F7F),
    .INIT_53(256'h0000000000000000FF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FF),
    .INIT_54(256'h7F0000FFFFFFFFFFFFFFFFFF7F7F7F7F7F7F7F7F7F00007F7F7F7F7F7F7F7F7F),
    .INIT_55(256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F),
    .INIT_56(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFF00007F7F7F7F7F),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h808080808080808098B8F0E0C080000000000000000000000000000000000000),
    .INIT_5C(256'h808080808080808000000000000080C0E0F0F0E0C08000000000000080808080),
    .INIT_5D(256'h000000000000000000FFFF000000000000000000000080C0E0F0B89880808080),
    .INIT_5E(256'h0000C0E06070381C0E0607030000000000000080C0C0E0E0E0FEFCF8F0E0C000),
    .INIT_5F(256'h000000000307060E1C387060E0C0000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h6070381C0C060703000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0307060E1C387060E0C0C0E06070381C0C06070300000000000000000000C0E0),
    .INIT_63(256'hE0C0800000000000000000000307060E1C387060E0C000000000000000000000),
    .INIT_64(256'h0E06070300000000000000000080C0E06070381C0E0607030307060E1C387060),
    .INIT_65(256'h1C387060E0C0C0E06070381C0C0607030307060C1C387060E0C0C0E06070381C),
    .INIT_66(256'hFCFCF8F0E0C08000000000006070787CFEFFFFFE7C787060000000000307060E),
    .INIT_67(256'h0307060E1C387060E0C0C0E06070381C0C0607030080C0E0F0F8FCFCC0C0C0C0),
    .INIT_68(256'h00010307060E1C387060E0C0000000000000C0F0F8F87C3C3C3C3C3C00000000),
    .INIT_69(256'h7060E0C0C0E06070381C0E060703010000000000000000000000000000000000),
    .INIT_6A(256'h00000000000000000000000000000000C0E06070381C0E0607030307060E1C38),
    .INIT_6B(256'h0000000000000000800000000000000000010307060E1C387060E0C080000000),
    .INIT_6C(256'hC0E06070381C0E0607030307060E1C387060E0C0C0E06070381C0E0607030100),
    .INIT_6D(256'h00010307060E1C387060E0C00000000000000000000000000000000000000080),
    .INIT_6E(256'h7060E0C0C0E06070381C0E060703010000000000000000800000000000000000),
    .INIT_6F(256'h00000000000000000000000000000080C0E06070381C0E0607030307060E1C38),
    .INIT_70(256'h0000000000000080800000000000000000010307060E1C387060E0C080000000),
    .INIT_71(256'hC0E06070381C0E0607030307060E1C387060E0C0C0E06070381C0E0607030100),
    .INIT_72(256'h0F0F0F0F1C38F8E00000000000000000E0F8381C0C0C0C0C1C38F8E0C0C0C0C0),
    .INIT_73(256'h00000000C0C0C0C0E0F8381C0C0C0C0C1C38F8E00000000000000000E0F8381C),
    .INIT_74(256'hE0F8381C0C0C0C0C1C38F8E0C0C0C0C000000000E0F8381C0C0C0C0C1C38F8E0),
    .INIT_75(256'hFCF8F8E0C0C0C0C000000000E0F8381C0F0F0F0F1C38F8E000000000C0C0C0C0),
    .INIT_76(256'h00000000E0F8F8FCFFFFFFFFFCF8F8E00000000000000000E0F8F8FCFCFCFCFC),
    .INIT_77(256'hFCFCFCFCFCF8F8E000000000C0C0C0C0E0F8F8FCFCFCFCFCFCF8F8E000000000),
    .INIT_78(256'h00000000C0C0C0C0E0F8F8FCFCFCFCFCFCF8F8E0C0C0C0C000000000E0F8F8FC),
    .INIT_79(256'hF8F0E0C080000000000000000000000000000000E0F8F8FCFFFFFFFFFCF8F8E0),
    .INIT_7A(256'hC0E0F0F8FCFCC0C00000000000000000008080000000000000000000C0C0FCFC),
    .INIT_7B(256'h000000000C1C3C7CFFFFFFFF7C3C1C0C00000000000000000000000000000080),
    .INIT_7C(256'hE080000000000000000000000000000000000000FFFF00000000000000000000),
    .INIT_7D(256'h0000000000000000000000003F7FE0C0808000000000000000000C0C1C1838F0),
    .INIT_7E(256'h1C1838F0E080000000000000000000000000000000000000E0F83C0C07070303),
    .INIT_7F(256'h00000000000000000000000000000000F0F83C0C070703030000000000000C0C),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_20480x16_sub_008192_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_Naddra[12]_addra_o ),
    .dia({open_n279,open_n280,open_n281,open_n282,open_n283,open_n284,open_n285,open_n286,dia[7:0]}),
    .wea(wea),
    .doa({open_n308,open_n309,open_n310,open_n311,open_n312,open_n313,open_n314,open_n315,inst_doa_i2_007,inst_doa_i2_006,inst_doa_i2_005,inst_doa_i2_004,inst_doa_i2_003,inst_doa_i2_002,inst_doa_i2_001,inst_doa_i2_000}));
  // address_offset=8192;data_offset=8;depth=4096;width=8;num_section=1;width_per_section=8;section_size=16;working_depth=4096;working_width=8;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h020202020000000000000000FF0000FF00000000000000000000000000000000),
    .INIT_01(256'h02020202FE0000FF00000000000000000000000000000000FF0000FE02020202),
    .INIT_02(256'h00000000000000000202020202020202FE0000FE020202020202020202020202),
    .INIT_03(256'h0202020202020202FE0000FE02020202020202020202020202020202FE0000FF),
    .INIT_04(256'h0303030303030303030303030000000000000000030303030000000000000000),
    .INIT_05(256'h0303030300000000000000000303030300000000000000000000000000000000),
    .INIT_06(256'h0303030303030303000000000000000000000000000000000303030303030303),
    .INIT_07(256'h0000000000000000030303030303030303030303030303030303030303030303),
    .INIT_08(256'h0303030303030303030303030303030303030303030303030303030303030303),
    .INIT_09(256'hFFFFFFFF03030303030303030000000000000000FFFFFFFF0000000000000000),
    .INIT_0A(256'h030303030000000000000000FFFFFFFF00000000000000000000000000000000),
    .INIT_0B(256'h03030303FFFFFFFF00000000000000000000000000000000FFFFFFFF03030303),
    .INIT_0C(256'h00000000000000000303030303030303FFFFFFFF030303030303030303030303),
    .INIT_0D(256'h0303030303030303FFFFFFFF03030303030303030303030303030303FFFFFFFF),
    .INIT_0E(256'h0100000101010100000101010202020000020202020000020202020000020202),
    .INIT_0F(256'h0000000003030300000303030300000303030300000303030101010000010101),
    .INIT_10(256'h0000000000CECE0000000000000000000000000000000000CE0000CE00000000),
    .INIT_11(256'h02020202020202020000000000000000CECECECE000000000000000000000000),
    .INIT_12(256'h020202020202020202FEFE020202020202020202020202020202020202020202),
    .INIT_13(256'hFF0000FF00000000000000000000000000000000FF0000FF0101010101010101),
    .INIT_14(256'h030303030303030303030303FFFFFFFF01010101010101010101010101010101),
    .INIT_15(256'h01010101FFFFFFFF0303030303030303030303030303030303FFFF0303030303),
    .INIT_16(256'h01010101010101010303030303030303FFFFFFFF030303030303030301010101),
    .INIT_17(256'h030303030303030303FFFF0303030303030303030101010101010101FFFFFFFF),
    .INIT_18(256'h0101010101010101010101010000000000000000000303030303030303030303),
    .INIT_19(256'h0000000003030303030303030303030000000000000000000000000000000000),
    .INIT_1A(256'h0000000000FFFF03030303030303030301010101010101010101010100000000),
    .INIT_1B(256'h00000000000000000000000000000000FFFFFFFF010101010101010100000000),
    .INIT_1C(256'h0101010101010101FFFFFFFF0000000000000000030303030303030303FFFF00),
    .INIT_1D(256'h0101010101010101010101010303030303030303030303030303030303030303),
    .INIT_1E(256'h01010101030303030303030303FFFF0303030303030303030101010101010101),
    .INIT_1F(256'h00000000FFFFFFFF01010101010101010101010101010101FFFFFFFF01010101),
    .INIT_20(256'h0000000000000000000000000000000000FFFF03030303030303030300000000),
    .INIT_21(256'h030303030303030303FFFF0000000000000000000101010101010101FFFFFFFF),
    .INIT_22(256'h0303030302020202020202020000000000000000030303030303030303030303),
    .INIT_23(256'h0000000003030303030303030303030300000000000000000000000000000000),
    .INIT_24(256'h00000000FF0303FF030303030303030302020202020202020303030300000000),
    .INIT_25(256'h00000000000000000000000000000000FFFFFFFF020202020202020200000000),
    .INIT_26(256'h0202020202020202FFFFFFFF00000000000000000303030303030303FF0303FF),
    .INIT_27(256'h0202020202020202020202020303030303030303030303030303030303030303),
    .INIT_28(256'h0202020202020202020202020303030303030303030303030202020202020202),
    .INIT_29(256'h03030303FF0303FF030303030303030303030303030303030303030302020202),
    .INIT_2A(256'h03030303030303030202020202020202FEFEFEFE020202020202020203030303),
    .INIT_2B(256'h0303030303030303FFFFFFFF02020202020202020202020202020202FFFFFFFF),
    .INIT_2C(256'hFFFFFFFF03030303030303030202020202020202FF0303FF0303030303030303),
    .INIT_2D(256'h030303030303030303030303FFFFFFFF02020202020202020202020202020202),
    .INIT_2E(256'h02020202FFFFFFFF03030303030303030303030303030303FF0303FF03030303),
    .INIT_2F(256'h03030303030303030303030303030303FFFFFFFF030303030303030302020202),
    .INIT_30(256'h0202020202020202FEFEFEFE02020202020202020303030303030303FF0000FF),
    .INIT_31(256'hFFFFFFFF02020202020202020000000000000000FF0000FF0303030303030303),
    .INIT_32(256'h030303030000000000000000FFFFFFFF03030303030303030000000000000000),
    .INIT_33(256'h03030303FF0303FF00000000000000000000000000000000FF0303FF03030303),
    .INIT_34(256'h00000000000000000303030303030303FFFFFFFF000000000000000003030303),
    .INIT_35(256'h0303030303030303FF0000FF00000000000000000202020202020202FFFFFFFF),
    .INIT_36(256'hFF0303FF02020202020202020303030303030303FFFFFFFF0202020202020202),
    .INIT_37(256'h000000000000000000000000FFFFFFFF00000000000000000303030303030303),
    .INIT_38(256'h030303030303020202020202020202020000000000000000FF0000FF00000000),
    .INIT_39(256'h0101010101010101020202020202020202020303030303030303030303030303),
    .INIT_3A(256'h0101010101010101FF0101FF0101010101010101010101010101010101010101),
    .INIT_3B(256'h02FFFF000000000000000000000000000000000000FFFF020202020202020202),
    .INIT_3C(256'hFFFFFFFFFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE0202020202020202),
    .INIT_3D(256'h02020202020202020202020202020202FFFFFFFFFFFFFFFFFF0000FFFFFFFFFF),
    .INIT_3E(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE0000FF000000000000000002020202),
    .INIT_3F(256'h0000000000000000FF0000FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE0000FE),
    .INIT_40(256'h0202020202020202020202020202020202020202020202020202020202020202),
    .INIT_41(256'h000000000202020202020202FE0000FF00000000000000000202020202020202),
    .INIT_42(256'hFEFEFEFEFE0000FE0202020202020202FEFEFEFEFEFEFEFEFE0000FF00000000),
    .INIT_43(256'hFEFEFEFEFEFEFEFE0202020202020202FE0000FEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_44(256'h0000000000000000FF0000FE02020202020202020000000000000000FF0000FE),
    .INIT_45(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_46(256'hFFFFFFFF0202020202020202FE0000FFFFFFFFFFFFFFFFFFFEFEFEFEFEFEFEFE),
    .INIT_47(256'hFEFEFEFEFE0000FE0202020202020202FEFEFEFEFEFEFEFEFE0000FFFFFFFFFF),
    .INIT_48(256'hFEFEFEFEFEFEFEFE0202020202020202FE0000FEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_49(256'hFFFFFFFFFFFFFFFFFF0000FE0202020202020202FFFFFFFFFFFFFFFFFF0000FE),
    .INIT_4A(256'h0302020202020202020202020202020202020202020202030000000000000000),
    .INIT_4B(256'h000000000000000000000000FF0000FEFEFEFEFEFEFEFEFE0000000000000000),
    .INIT_4C(256'hFEFEFEFEFEFEFEFFFFFFFFFFFFFFFFFFFEFEFEFEFEFEFEFEFE0000FF00000000),
    .INIT_4D(256'h0202020202020202FFFFFFFFFFFFFFFFFFFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_4E(256'h0202020202020202FE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FE),
    .INIT_4F(256'hFFFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFFFFFFFFFFF),
    .INIT_50(256'hFFFFFFFFFFFFFFFFFFFFFFFFFF0000FEFEFEFEFEFEFEFEFEFFFFFFFFFFFFFFFF),
    .INIT_51(256'h02020202020202020202020202020202FEFEFEFEFEFEFEFEFE0000FFFFFFFFFF),
    .INIT_52(256'h0000000000000000FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE02020202),
    .INIT_53(256'h0000000000000000FF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FF),
    .INIT_54(256'hFE0000FFFFFFFFFFFFFFFFFFFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_55(256'hFEFEFEFEFEFEFEFEFEFEFEFEFE0000FEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_56(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFF0000FEFEFEFEFE),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0101010101010101191D0F070301000000000000000000000000000000000000),
    .INIT_5C(256'h0101010101010101000000000003030100FFFF00010303000000000001010101),
    .INIT_5D(256'h000000000003070E1C3F3F1C0E0703000000000000000103070F1D1901010101),
    .INIT_5E(256'h0000000000000000000000000000000000007E7F7F7F0301011F0F0703010000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000307060E1C387060E0C0C0E06070381C0E060703000000000000),
    .INIT_61(256'h060E1C383060E0C0C0E06070381C0E0607030307060E1C383060E0C000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000307),
    .INIT_63(256'h07030307060E1C383060E0C0C0E06070381C0E06070300000000000000000000),
    .INIT_64(256'h7060E0C0C0E06030381C0E0607030307060E1C387060E0C0C0E06070381C0E06),
    .INIT_65(256'h381C0E06070301000000000000000000000000000000000000010307060E1C38),
    .INIT_66(256'h3F3F1F0F0703010000000000060E1E3E7FFFFF7F3E1E0E0600000000C0E06070),
    .INIT_67(256'hC0E06070381C0E0607030307060E1C383060E0C0000103070F1F3F3F03030303),
    .INIT_68(256'h000000000000000000000001000002060E1E3F7F7F3F1E0E0602000000000000),
    .INIT_69(256'h0000000101000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h1C387060E0C08000000000000000000001000000000000000000000000000000),
    .INIT_6B(256'h00000000000000000307060E1C387060E0C0800000000000000000010307060E),
    .INIT_6C(256'h0307060E1C387060E0C0800000000000000000010307060E1C387060E0C08000),
    .INIT_6D(256'h0080C0E06070381C0E06070300000000000000000080C0E06070381C0E060703),
    .INIT_6E(256'h0E06070301000000000000000080C0E06070381C0E0607030000000000000000),
    .INIT_6F(256'h1C387060E0C0C0E06070381C0E06070301000000000000000080C0E06070381C),
    .INIT_70(256'h6070381C0E0607030307060E1C387060E0C0C0E06070381C0E0607030307060E),
    .INIT_71(256'h0307060E1C387060E0C0C0E06070381C0E0607030307060E1C387060E0C0C0E0),
    .INIT_72(256'h30303030381C1F070000000000000000071F1C3830303030381C1F0703030303),
    .INIT_73(256'h0000000003030303071F1C3830303030381C1F070000000000000000071F1C38),
    .INIT_74(256'h071F1C3830303030381C1F070303030300000000071F1C38F0F0F0F0381C1F07),
    .INIT_75(256'h3F1F1F070303030300000000071F1C38F0F0F0F0381C1F070000000003030303),
    .INIT_76(256'h00000000071F1F3F3F3F3F3F3F1F1F070000000000000000071F1F3F3F3F3F3F),
    .INIT_77(256'hFFFFFFFF3F1F1F070000000003030303071F1F3F3F3F3F3F3F1F1F0700000000),
    .INIT_78(256'h0000000003030303071F1F3F3F3F3F3F3F1F1F070303030300000000071F1F3F),
    .INIT_79(256'h1F0F070301000000000000000000000000000000071F1F3FFFFFFFFF3F1F1F07),
    .INIT_7A(256'h03070F1F3F3F03030000000030383C3EFFFFFFFF3E3C38300000000003033F3F),
    .INIT_7B(256'h0000000000000000000101000000000000000000000000000000000000000001),
    .INIT_7C(256'hFFFF000000000000000000000000C0C0E060703C1F0700000000000000000000),
    .INIT_7D(256'h000000000000000000000000F0F81C0C07070303000000000000000000000000),
    .INIT_7E(256'h000000003F7FE0C080800000000000000000C0C0E060703C1F07000000000000),
    .INIT_7F(256'h80800000000000000000000000000000FFFF0000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_20480x16_sub_008192_008 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_Naddra[12]_addra_o ),
    .dia({open_n336,open_n337,open_n338,open_n339,open_n340,open_n341,open_n342,open_n343,dia[15:8]}),
    .wea(wea),
    .doa({open_n365,open_n366,open_n367,open_n368,open_n369,open_n370,open_n371,open_n372,inst_doa_i2_015,inst_doa_i2_014,inst_doa_i2_013,inst_doa_i2_012,inst_doa_i2_011,inst_doa_i2_010,inst_doa_i2_009,inst_doa_i2_008}));
  // address_offset=12288;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=16;working_depth=4096;working_width=8;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h00000000000000000000FFFF00000000000000000000000000000000FFFF0000),
    .INIT_01(256'hC0E07F3F00000000000000000000000000000000000080E0F038181C0C0C0000),
    .INIT_02(256'h0C0C000000000000030307070C3CF8E000000000000000000000000000008080),
    .INIT_03(256'h030307070C3CF8F000000000000000000000000000000000000080E0F038181C),
    .INIT_04(256'h808080000000000000000000000000000000FFFF000000000000000000000000),
    .INIT_05(256'hC0C0C0C0C0C08000000000808080C0E060703C1C000000000080C0F03C3CF0C0),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h000000000000000000000080C0F03C3CF0C08000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000080C0F03C3CF0C0800000000000000000000000),
    .INIT_09(256'h000000000080C0F03C3CF0C08000000000000000000000000000000000000000),
    .INIT_0A(256'hC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0E060703C1C000000000000000000000000),
    .INIT_0B(256'h800000000080C0C0C0C0C0C000001C3C7060E0C0C0C0C0C0C0C0C0C0C0C0C0C0),
    .INIT_0C(256'hC0C0800000000080C0C0C0C0C0C0C0C0C0C0C0E060703C1CC0C0C0C0C0C0C0C0),
    .INIT_0D(256'hC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C000001C3C7060E0C0C0C0C0C0C0C0C0C0),
    .INIT_0E(256'h0080C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0800000000080),
    .INIT_0F(256'h0000000000000080C0F03C3CF0C080000000000000001C3C7060E0C080000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'hC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C000000000000000000000000000000000),
    .INIT_13(256'h0C0C0C0C0C0C0C0C3030303030303030303030303030303030303030C0C0C0C0),
    .INIT_14(256'h03030303030303030303030303030303030303030C0C0C0C0C0C0C0C0C0C0C0C),
    .INIT_15(256'hFCFCF0C000000000000000000303070F3EFCF0C00000C0F0FC3E0F0703030303),
    .INIT_16(256'h0000000000000000000000008080C0C0E0E07070383C1F0F000000000000C0F0),
    .INIT_17(256'h3FFFFFFFFFFFFFFFFF3F0F03030303030F1F3C387070E0E0C0C0808000000000),
    .INIT_18(256'hE0E0F0F0F8F8FFFF000000000000C0F0FCFCF0C000000000000000000303030F),
    .INIT_19(256'hFFFFF8F8F0F0E0E0C0C08080000000000000000000000000000000008080C0C0),
    .INIT_1A(256'h0000000000000000FFFF0000000000000000000000000000000000000000FFFF),
    .INIT_1B(256'h000000000000000000000000000000000000FFFF000000000000000000000000),
    .INIT_1C(256'h000000000000FFFF0000000000000000000000000000000000000000FFFF0000),
    .INIT_1D(256'h00000000000000000000000000000000FFFF0000000000000000000000000000),
    .INIT_1E(256'h00000000FFFF0000000000000000000000000000000000000000FFFF00000000),
    .INIT_1F(256'h0000000000000000000000000000FFFF00000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000F1F3830E0E0C0C000000000FFFF000000000000),
    .INIT_21(256'h00000000000080E0F038181C0C0C000000000000C0C0E0E030381F0F00000000),
    .INIT_22(256'h000000000000000000000C0C1C1838F0E0800000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h000000000000000000000000000000000000000000000000FEF8C00000000000),
    .INIT_26(256'h00000000000000000000000000000000FFFCF8F0E0C080000000000000000000),
    .INIT_27(256'hFFFFFFFFFFFFFFFFFFFEFCF8F0F0E0C080000000000000000000000000000000),
    .INIT_28(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F0F03FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_29(256'hFFFFFFFFFFFF3F1F0F070301FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2A(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2B(256'hFFFFFFFFFF7F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F1F07010000),
    .INIT_2C(256'hC080800000000000FFFFFFFFFFFFFFFFFFFFFFFFFF7F3F1F0F070301FFFFFFFF),
    .INIT_2D(256'h00000000000080C0E0F0F0E0C0800000000000000000000000F8F8F0F0E0E0C0),
    .INIT_2E(256'h000000000000000000000000FF3F1F0703010000000000000000000000000000),
    .INIT_2F(256'h00000000FF7F7F3F1F1F0F0F070703030101000000000000FFFFFF7F0F030000),
    .INIT_30(256'h3F3F1F1F1F0F0F0F0707070303030101FFFFFFFFFFFFFF7F3F1F0F0301000000),
    .INIT_31(256'hFFFFFFFCF8E0C080FFFFFFFFFFFFFFFFFFFFFF7F3F1F0F0F07030301FF7F7F7F),
    .INIT_32(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF0C0000000FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_33(256'hF8F0E0C08000000000000000FFFFFFFFFFFFFFFEFEFCF8F8F0F0E0E0C0808000),
    .INIT_34(256'h00000000FFFEFEFEFCFCF8F8F8F0F0E0E0E0C0C080808000FFFFFFFFFFFFFEFC),
    .INIT_35(256'hF0E0C0800000000080C0E0F0F8FCFEFFFFFFFFFFFFFFFEF8E080000000000000),
    .INIT_36(256'hF0F8F800000000000103070F1F3F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFCF8),
    .INIT_37(256'h0000002060E0E0E0E0E0E0E0E0E0E0602000000000000000008080C0C0E0E0F0),
    .INIT_38(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_39(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF030F7FFFFFFFFFFF),
    .INIT_3A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000001030F1F3F7FFFFFFF),
    .INIT_3B(256'h0000000000000000010303070F0F1F3F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_3C(256'h0000000000000000000000000000000000C0F8FE000000000000000000000000),
    .INIT_3D(256'h000000000080C0E0F0F8FCFE0000000000000000000000000000000000000000),
    .INIT_3E(256'hFFFFFFFF00000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h000000000080800000000000000000000000000000000000000080E0F8FEFFFF),
    .INIT_40(256'hC0C08080000000000000000000000000000000000080C0E0F0F8FCFE00000000),
    .INIT_41(256'h0000000000000080C0E0E0C08000000000000000FFFFFEFEFCFCF8F8F0F0E0E0),
    .INIT_42(256'hFFFFFFFFFFFFFFFFFFFFFFFF80C0E0F8FCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_43(256'hF0F8FCFF008080C0E0E0F0F0F8F8FCFEFEFFFFFFFFFFFFFF000000C0F0FCFFFF),
    .INIT_44(256'hC0C0E0E0E0F0F0F8F8F8FCFCFEFEFEFF0000000000000000000000000080C0E0),
    .INIT_45(256'h00000103071F3FFF000000000000000000000080C0E0F0F0F8FCFEFF00808080),
    .INIT_46(256'h0000000000000000000000000000030F7FFFFFFF000000000000000000000000),
    .INIT_47(256'h030F1F3F7FFFFFFFFFFFFFFF0000000000000101030307070F0F1F1F3F7F7FFF),
    .INIT_48(256'hFFFFFFFF01010303030707070F0F0F1F1F1F3F3F7F7F7FFF0000000000000001),
    .INIT_49(256'h0F1F3F7FFFFFFFFF7F3F1F0F0703010000000000000001071F7FFFFFFFFFFFFF),
    .INIT_4A(256'hF8F8FCFCFEFEFFFFFEFCF8F0E0C0800000000000000000000000000000010307),
    .INIT_4B(256'h03070F1F3F7FFFFFFFFFFFFFFFFF7F3F1F0F0703000000008080C0C0E0E0F0F0),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'hC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C000000000000000000000000000000000),
    .INIT_4F(256'hFCFCFCFCFCFCFCFCF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0C0C0C0C0),
    .INIT_50(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFCFCFCFCFCFCFCFCFCFCFC),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'hC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C000000000000000000000000000000000),
    .INIT_54(256'hFCFCFCFCFCFCFCFC0000F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F00000C0C0),
    .INIT_55(256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FCFCFCFCFCFCFCFCFCFC),
    .INIT_56(256'h0F0F0F0F0F0F0F0F0F0F0F0F0303030303030303030303030303030303030303),
    .INIT_57(256'hFFFFFFFF3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F0F0F0F0F0F0F0F0F),
    .INIT_58(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_59(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5B(256'h0F0F0F0F0F0F0F0F0F0F0F0F0000010101010101010101010101010101010101),
    .INIT_5C(256'hFFFFFFFF00003F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F00000F0F0F0F0F0F),
    .INIT_5D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5E(256'hFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFF),
    .INIT_5F(256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFF),
    .INIT_60(256'h000000000000000000000000FFFF000000000000000000000000000000000000),
    .INIT_61(256'h00000000FFFFFFFFFFFF0000000000000000000000000000FFFFFFFF00000000),
    .INIT_62(256'hFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFFFFFF0000000000000000),
    .INIT_63(256'hFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000FFFFFFFF),
    .INIT_64(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_65(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000),
    .INIT_66(256'h03030303030303030303030303030303030303030303FFFFFFFFFFFFFFFFFFFF),
    .INIT_67(256'h00000000000000000000000000000000FFFF0303030303030303030303030303),
    .INIT_68(256'h000000000000FFFF000000000000000000000000000000000000FFFFFFFF0000),
    .INIT_69(256'h0303030303030303030303030303030303030303FFFF00000000000000000000),
    .INIT_6A(256'h000000000000000000000000FCFC000000000000000000000000000000000000),
    .INIT_6B(256'h00000000FCFCFCFCFCFC0000000000000000000000000000FCFCFCFC00000000),
    .INIT_6C(256'hFCFCFCFCFCFC00000000000000000000FCFCFCFCFCFCFCFC0000000000000000),
    .INIT_6D(256'hFCFC000000000000FCFCFCFCFCFCFCFCFCFCFCFC0000000000000000FCFCFCFC),
    .INIT_6E(256'hFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC00000000FCFCFCFCFCFCFCFCFCFCFCFC),
    .INIT_6F(256'hFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC0000),
    .INIT_70(256'h03030303FFFF03030303030303030303030303030303FFFFFCFCFCFCFCFCFCFC),
    .INIT_71(256'h0000000000000000000000000000FFFFFFFF0303030303030303030303030303),
    .INIT_72(256'h030303030303FFFF030303030303030303030303030303030303FFFFFFFF0000),
    .INIT_73(256'h0000000000000000000000000000000000000000FFFF03030303030303030303),
    .INIT_74(256'h0000000000000000FFFFFFFF000000000000000000000000000000000000FFFF),
    .INIT_75(256'hFFFFFFFF0000000000000000000000000000FFFFFFFFFFFF0000000000000000),
    .INIT_76(256'h000000000000FFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
    .INIT_77(256'hFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFF00000000),
    .INIT_78(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF),
    .INIT_79(256'hFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_7A(256'h000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFF),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000FCFCFCFC000000000000000000000000000000000000FCFC),
    .INIT_7F(256'hFCFCFCFC0000000000000000000000000000FCFCFCFCFCFC0000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_20480x16_sub_012288_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_addra[12]_addra[_o ),
    .dia({open_n393,open_n394,open_n395,open_n396,open_n397,open_n398,open_n399,open_n400,dia[7:0]}),
    .wea(wea),
    .doa({open_n422,open_n423,open_n424,open_n425,open_n426,open_n427,open_n428,open_n429,inst_doa_i3_007,inst_doa_i3_006,inst_doa_i3_005,inst_doa_i3_004,inst_doa_i3_003,inst_doa_i3_002,inst_doa_i3_001,inst_doa_i3_000}));
  // address_offset=12288;data_offset=8;depth=4096;width=8;num_section=1;width_per_section=8;section_size=16;working_depth=4096;working_width=8;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h00000000000000000000071F3C7060E0C0C0000000000000000000003F7FE0C0),
    .INIT_01(256'h0C1CF8F0000000000000000000000000000000000000FFFF0000000000000000),
    .INIT_02(256'h0000000000000000000000000000071F3C7060E0C0C000000000000003030707),
    .INIT_03(256'h000000000000FFFF00000000000000000000000000008080C0E07F3F00000000),
    .INIT_04(256'h01010307060E3C380000000000008080C0E07F3F000000000000000000000000),
    .INIT_05(256'h000000000001030F3C3C0F030101010000000000030303030303010000000001),
    .INIT_06(256'h03030303030303030303030303030303030303030303030303030307060E3C38),
    .INIT_07(256'h060E3C3803030303030303030100000000010303030303030000383C0E060703),
    .INIT_08(256'h0E06070303030303030303030303010000000001030303030303030303030307),
    .INIT_09(256'h030303030303010000000001030303030303030303030303030303030000383C),
    .INIT_0A(256'h0000000000000000000000000000000000000000030303030303030303030303),
    .INIT_0B(256'h030F3C3C0F030100000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0001030F3C3C0F03010000000000000000000000000000000000000000000001),
    .INIT_0D(256'h0100000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0F03010000000000000000000000000000000000000000000001030F3C3C0F03),
    .INIT_0F(256'h0000383C0E0607030100000000010303030303030000000000000001030F3C3C),
    .INIT_10(256'h303030303030303030303030C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0),
    .INIT_11(256'h030303030C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C3030303030303030),
    .INIT_12(256'h0000000000000000000000000000000003030303030303030303030303030303),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000030F3F7CF0E0C0C0C0C0000000000000030F3F3F0F030000000000000000),
    .INIT_16(256'h00000000000000000000030307070F0F1C1C383870F0E0C0C0C0E0F07C3F0F03),
    .INIT_17(256'h0000030F3F3F0F030000000000000000C0E0F07038381C1C0F0F070703030000),
    .INIT_18(256'h1F1F3F3F7F7FFFFFC0C0C0F0FCFFFFFFFFFFFFFFFFFCF0C0C0C0C0C000000000),
    .INIT_19(256'hFFFF7F7F3F3F1F1F0F0F07070303000000000000000000000000030307070F0F),
    .INIT_1A(256'h0000000000000000FFFF0000000000000000000000000000000000000000FFFF),
    .INIT_1B(256'h000000000000000000000000000000000000FFFF000000000000000000000000),
    .INIT_1C(256'h000000000000FFFF0000000000000000000000000000000000000000FFFF0000),
    .INIT_1D(256'h00000000000000000000000000000000FFFF0000000000000000000000000000),
    .INIT_1E(256'h00000000FFFF0000000000000000000000000000000000000000FFFF00000000),
    .INIT_1F(256'h0000000000000000000000000000FFFF00000000000000000000000000000000),
    .INIT_20(256'hC0C000000000C0C0E060703C1E0603030101000000000000FFFF000000000000),
    .INIT_21(256'h0C0C1E1E3373E1C1000000000000000000000000000001010303061E3C7060E0),
    .INIT_22(256'h00000000000000000000000000000000C1E173331E1E0C0C0000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h000000000000000000000000FFFCF8E0C0800000000000000000000000000000),
    .INIT_25(256'h00000000FFFEFEFCF8F8F0F0E0E0C0C08080000000000000FFFFFFFEF0C00000),
    .INIT_26(256'hFCFCF8F8F8F0F0F0E0E0E0C0C0C08080FFFFFFFFFFFFFFFEFCF8F0C080000000),
    .INIT_27(256'hFFFFFF3F1F070301FFFFFFFFFFFFFFFFFFFFFFFEFCF8F0F0E0C0C080FFFEFEFE),
    .INIT_28(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF3F0F03000000FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_29(256'h1F0F07030100000000000000FFFFFFFFFFFFFF7F7F3F1F1F0F0F070703010100),
    .INIT_2A(256'h00000000FF7F7F7F3F3F1F1F1F0F0F070707030301010100FFFFFFFFFFFF7F3F),
    .INIT_2B(256'h0F070301000000000103070F1F3F7FFFFFFFFFFFFFFF7F1F0701000000000000),
    .INIT_2C(256'h0301010000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFEFCF8F0E0C080FF7F3F1F),
    .INIT_2D(256'h000000040607070707070707070707060400000000000000001F1F0F0F070703),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000007F1F030000000000),
    .INIT_30(256'h00000000000000000000000000000000FF3F1F0F070301000000000000000000),
    .INIT_31(256'hFFFFFFFFFFFFFFFFFF7F3F1F0F0F070301000000000000000000000000000000),
    .INIT_32(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF0C0FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_33(256'hFFFFFFFFFFFFFCF8F0E0C080FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_34(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_35(256'hFFFFFFFFFFFEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF8E0800000),
    .INIT_36(256'h0F1F1F000000000080C0E0F0F8FCFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_37(256'h0000000000000103070F0F07030100000000000000000000000101030307070F),
    .INIT_38(256'hFFFFFFFFFFFFFFFFFFFFFFFF0103071F3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_39(256'h0F1F3FFF0001010307070F0F1F1F3F7F7FFFFFFFFFFFFFFF000000030F3FFFFF),
    .INIT_3A(256'h03030707070F0F1F1F1F3F3F7F7F7FFF00000000000000000000000000010307),
    .INIT_3B(256'h000080C0E0F8FCFF00000000000000000000000103070F0F1F3F7FFF00010101),
    .INIT_3C(256'h0000000000000000000000000000C0F0FEFFFFFF000000000000000000000000),
    .INIT_3D(256'hC0F0F8FCFEFFFFFFFFFFFFFF0000000000008080C0C0E0E0F0F0F8F8FCFEFEFF),
    .INIT_3E(256'hFFFFFFFF8080C0C0C0E0E0E0F0F0F0F8F8F8FCFCFEFEFEFF0000000000000080),
    .INIT_3F(256'hF0F8FCFEFFFFFFFFFEFCF8F0E0C0800000000000000080E0F8FEFFFFFFFFFFFF),
    .INIT_40(256'h0303010100000000000000000000000000000000000103070F1F3F7F0080C0E0),
    .INIT_41(256'hC0E0F0F8FCFEFFFFFFFFFFFFFFFFFEFCF8F0E0C0FFFF7F7F3F3F1F1F0F0F0707),
    .INIT_42(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_43(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0F0FEFFFFFFFFFF),
    .INIT_44(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000080C0F0F8FCFEFFFFFF),
    .INIT_45(256'h000000000000000080C0C0E0F0F0F8FCFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_46(256'h0000000000000000000000000000000000031F7F000000000000000000000000),
    .INIT_47(256'h00000000000103070F1F3F7F0000000000000000000000000000000000000000),
    .INIT_48(256'hFFFFFFFF00000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h000000000001010000000000000000000000000000000000000001071F7FFFFF),
    .INIT_4A(256'h1F1F3F3F7F7FFFFF7F3F1F0F0703010000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000001030707030100000000000000000000000101030307070F0F),
    .INIT_4C(256'hF0F0F0F0F0F0F0F0F0F0F0F0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0),
    .INIT_4D(256'hFFFFFFFFFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF0F0F0F0F0F0F0F0),
    .INIT_4E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_4F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_50(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_51(256'hF0F0F0F0F0F0F0F0F0F0F0F00000808080808080808080808080808080808080),
    .INIT_52(256'hFFFFFFFF0000FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC0000F0F0F0F0F0F0),
    .INIT_53(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_54(256'hFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFF),
    .INIT_55(256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFF),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0303030303030303030303030303030300000000000000000000000000000000),
    .INIT_59(256'h3F3F3F3F3F3F3F3F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F03030303),
    .INIT_5A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3F3F3F3F3F3F3F3F3F3F3F3F),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0303030303030303030303030303030300000000000000000000000000000000),
    .INIT_5E(256'h3F3F3F3F3F3F3F3F00000F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F00000303),
    .INIT_5F(256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00003F3F3F3F3F3F3F3F3F3F),
    .INIT_60(256'h000000000000000000000000FFFF000000000000000000000000000000000000),
    .INIT_61(256'h00000000FFFFFFFFFFFF0000000000000000000000000000FFFFFFFF00000000),
    .INIT_62(256'hFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFFFFFF0000000000000000),
    .INIT_63(256'hFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000FFFFFFFF),
    .INIT_64(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_65(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000),
    .INIT_66(256'h00000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFF),
    .INIT_67(256'hC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0FFFF0000000000000000000000000000),
    .INIT_68(256'h000000000000FFFFC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0FFFFFFFFC0C0),
    .INIT_69(256'hC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0FFFF00000000000000000000),
    .INIT_6A(256'h000000000000000000000000FFFF000000000000000000000000000000000000),
    .INIT_6B(256'h00000000FFFFFFFFFFFF0000000000000000000000000000FFFFFFFF00000000),
    .INIT_6C(256'hFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFFFFFF0000000000000000),
    .INIT_6D(256'hFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000FFFFFFFF),
    .INIT_6E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000),
    .INIT_70(256'hC0C0C0C0FFFF00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFF),
    .INIT_71(256'hC0C0C0C0C0C0C0C0C0C0C0C0C0C0FFFFFFFFC0C0C0C0C0C0C0C0C0C0C0C0C0C0),
    .INIT_72(256'hC0C0C0C0C0C0FFFFC0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0FFFFFFFFC0C0),
    .INIT_73(256'h0000000000000000000000000000000000000000FFFFC0C0C0C0C0C0C0C0C0C0),
    .INIT_74(256'h0000000000000000FFFFFFFF000000000000000000000000000000000000FFFF),
    .INIT_75(256'hFFFFFFFF0000000000000000000000000000FFFFFFFFFFFF0000000000000000),
    .INIT_76(256'h000000000000FFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
    .INIT_77(256'hFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFF00000000),
    .INIT_78(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF),
    .INIT_79(256'hFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_7A(256'h000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFF),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000FFFFFFFF000000000000000000000000000000000000FFFF),
    .INIT_7F(256'hFFFFFFFF0000000000000000000000000000FFFFFFFFFFFF0000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_20480x16_sub_012288_008 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_addra[12]_addra[_o ),
    .dia({open_n450,open_n451,open_n452,open_n453,open_n454,open_n455,open_n456,open_n457,dia[15:8]}),
    .wea(wea),
    .doa({open_n479,open_n480,open_n481,open_n482,open_n483,open_n484,open_n485,open_n486,inst_doa_i3_015,inst_doa_i3_014,inst_doa_i3_013,inst_doa_i3_012,inst_doa_i3_011,inst_doa_i3_010,inst_doa_i3_009,inst_doa_i3_008}));
  // address_offset=16384;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=16;working_depth=4096;working_width=8;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h000000000000FCFCFCFCFCFCFCFCFCFC000000000000000000000000FCFCFCFC),
    .INIT_01(256'hFCFCFCFCFCFCFCFC0000000000000000FCFCFCFCFCFCFCFCFCFCFCFC00000000),
    .INIT_02(256'h00000000FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC000000000000FCFCFCFCFCFC),
    .INIT_03(256'hFCFCFCFCFCFCFCFCFCFCFCFC0000FCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC),
    .INIT_04(256'h000000000000000000000000000000000000000000000000FCFCFCFCFCFCFCFC),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'hFEFEFEFEFCFCF8F8F0C00000FFFFFFFFFFFFFFFEFEFEFEFEFCFCF8F8F0C00000),
    .INIT_09(256'hFFFFFF0F0000C0F0F8F8FCFCFEFEFEFEFEFFFFFFFFFFFFFF0000C0F0F8F8FCFC),
    .INIT_0A(256'hFFFFFFFEFEFEFEFCFCFCF8F0E0C000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFF0000C0E0F0F8FCFCFCFEFEFEFEFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0F0FFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFEFEFEFEFCFCF8F8F0C000000000C0F0F8F8FCFCFEFEFEFEFCFCF8F8F0C00000),
    .INIT_0E(256'hF0C000000000C0F0F8F8FCFCFEFEFEFEFEFFFFFFFFFFFF0F0000C0F0F8F8FCFC),
    .INIT_0F(256'hFFFFFFFFFFFF7F7F7F3F3F1F1F0F07030FFFFFFFFFFFFFFEFEFEFEFEFCFCF8F8),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFEFEFCF8F0C000000000C0F0F8FCFEFEFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFF3F3FFFFFFFFFFFFFFFFFFF03070F1F1F3F3F7F7F7FFFFF),
    .INIT_12(256'h000000000000010103030F3F0000000000000000000000000000000000000000),
    .INIT_13(256'h000000003F0F0303010100000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000010103030F3F3F0F030301010000000000000000010103030F3F00000000),
    .INIT_16(256'h0000000000000000000000000000010103030F3F000000000000000000000000),
    .INIT_17(256'h0000000000000000000000003F0F030301010000000000000000000000000000),
    .INIT_18(256'h03030F3F00000000000000000000000000000000000000003F0F030301010000),
    .INIT_19(256'h010100000000000000000000000000003F0F0303010100000000000000000101),
    .INIT_1A(256'h0000010103030F3F0000000000000000000000000000010103030F3F3F0F0303),
    .INIT_1B(256'h3F0F030301010000000000000000010103030F3F3F0F03030101000000000000),
    .INIT_1C(256'h000000000000FFFF0000000000000000FFFF0000000000000000FFFF00000000),
    .INIT_1D(256'h0000000000000000FFFF0000000000000000FFFF0000000000000000FFFF0000),
    .INIT_1E(256'hFFFFF0F0F0F0F0F0F0F0FFFF0000000000000000FFFFC0C0C0C0C0C0C0C0FFFF),
    .INIT_1F(256'hFFFFFFFF0000000000000000FFFFFCFCFCFCFCFCFCFCFFFF0000000000000000),
    .INIT_20(256'h00000000FFFF0000000000000000FFFF0000000000000000FFFFFFFFFFFFFFFF),
    .INIT_21(256'h000000000000FFFF0000000000000000FFFF0000000000000000FFFF00000000),
    .INIT_22(256'h0000000000000000FFFF0000000000000000FFFF0000000000000000FFFF0000),
    .INIT_23(256'hFFFFC0C0C0C0C0C0C0C0FFFF0000000000000000FFFF0000000000000000FFFF),
    .INIT_24(256'hFCFCFFFF0000000000000000FFFFF0F0F0F0F0F0F0F0FFFF0000000000000000),
    .INIT_25(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000FFFFFCFCFCFCFCFC),
    .INIT_26(256'h303030303030F0F00000000000000000F0F03030303030303030F0F000000000),
    .INIT_27(256'h0000000000000000F0F03030303030303030F0F00000000000000000F0F03030),
    .INIT_28(256'hF0F03030303030303030F0F00000000000000000F0F03030303030303030F0F0),
    .INIT_29(256'h000000000000000000000000F0F0F0F0F0F0F0F0F0F0F0F00000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h3F3F3F3F000000000000000000000000000000003F3F3F3F0000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h000000003F3F3F3F000000000000000000000000000000000000000000000000),
    .INIT_34(256'h000000000000000000000000000000003F3F3F3F000000000000000000000000),
    .INIT_35(256'h3F3F3F3F3F3F00000000000000000000000000003F3F3F3F3F3F000000000000),
    .INIT_36(256'h3F3F3F3F00000000000000003F3F3F3F3F3F00003F3F3F3F0000000000000000),
    .INIT_37(256'h000000003F3F3F3F3F3F00000000000000000000000000003F3F3F3F3F3F0000),
    .INIT_38(256'h3F3F00003F3F3F3F00000000000000003F3F3F3F3F3F00000000000000000000),
    .INIT_39(256'h00000000000000003F3F3F3F3F3F00003F3F3F3F00000000000000003F3F3F3F),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h3F3F3F3F000000000000000000000000000000003F3F3F3F0000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h000000003F3F3F3F000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h000000000000000000000000000000003F3F3F3F000000000000000000000000),
    .INIT_3F(256'h3F3F3F3F3F3F00000000000000000000000000003F3F3F3F3F3F000000000000),
    .INIT_40(256'h3F3F3F3F00000000000000003F3F3F3F3F3F00003F3F3F3F0000000000000000),
    .INIT_41(256'h000000003F3F3F3F3F3F00000000000000000000000000003F3F3F3F3F3F0000),
    .INIT_42(256'h3F3F00003F3F3F3F00000000000000003F3F3F3F3F3F00000000000000000000),
    .INIT_43(256'h00000000000000003F3F3F3F3F3F00003F3F3F3F00000000000000003F3F3F3F),
    .INIT_44(256'h00000000000000000000000000003F3F3F3F0000000000000000000000000000),
    .INIT_45(256'h3F3F3F3F00003F3F3F3F000000000000000000003F3F3F3F00003F3F3F3F0000),
    .INIT_46(256'h3F3F000000000000000000000000000000003F3F3F3F00000000000000000000),
    .INIT_47(256'h000000003F3F3F3F00003F3F3F3F000000000000000000000000000000003F3F),
    .INIT_48(256'h00003F3F3F3F000000000000000000003F3F3F3F00003F3F3F3F000000000000),
    .INIT_49(256'h3F3F3F3F3F3F00000000000000003F3F3F3F00003F3F3F3F3F3F000000000000),
    .INIT_4A(256'h3F3F3F3F00003F3F3F3F00003F3F3F3F3F3F00003F3F3F3F00003F3F3F3F0000),
    .INIT_4B(256'h3F3F00003F3F3F3F3F3F00000000000000003F3F3F3F00003F3F3F3F3F3F0000),
    .INIT_4C(256'h3F3F00003F3F3F3F00003F3F3F3F00003F3F3F3F3F3F00000000000000003F3F),
    .INIT_4D(256'h00003F3F3F3F00003F3F3F3F3F3F00003F3F3F3F00003F3F3F3F00003F3F3F3F),
    .INIT_4E(256'h00000000000000000000000000003F3F3F3F0000000000000000000000000000),
    .INIT_4F(256'h3F3F3F3F00003F3F3F3F000000000000000000003F3F3F3F00003F3F3F3F0000),
    .INIT_50(256'h3F3F000000000000000000000000000000003F3F3F3F00000000000000000000),
    .INIT_51(256'h000000003F3F3F3F00003F3F3F3F000000000000000000000000000000003F3F),
    .INIT_52(256'h00003F3F3F3F000000000000000000003F3F3F3F00003F3F3F3F000000000000),
    .INIT_53(256'h3F3F3F3F3F3F00000000000000003F3F3F3F00003F3F3F3F3F3F000000000000),
    .INIT_54(256'h3F3F3F3F00003F3F3F3F00003F3F3F3F3F3F00003F3F3F3F00003F3F3F3F0000),
    .INIT_55(256'h3F3F00003F3F3F3F3F3F00000000000000003F3F3F3F00003F3F3F3F3F3F0000),
    .INIT_56(256'h3F3F00003F3F3F3F00003F3F3F3F00003F3F3F3F3F3F00000000000000003F3F),
    .INIT_57(256'h00003F3F3F3F00003F3F3F3F3F3F00003F3F3F3F00003F3F3F3F00003F3F3F3F),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'hFFFFFFFF0000000000000000000000000000FFFFFFFFFFFF0000000000000000),
    .INIT_5A(256'h000000000000000000000000000000000000000000000000000000000000FFFF),
    .INIT_5B(256'h0000FFFFFFFFFFFF000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000FFFFFFFFFFFF000000000000000000000000),
    .INIT_5D(256'hFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFF000000000000),
    .INIT_5E(256'hFFFFFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFF),
    .INIT_5F(256'h0000FFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFF),
    .INIT_60(256'hFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFFFFFF00000000000000000000),
    .INIT_61(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'hFFFFFFFF0000000000000000000000000000FFFFFFFFFFFF0000000000000000),
    .INIT_64(256'h000000000000000000000000000000000000000000000000000000000000FFFF),
    .INIT_65(256'h0000FFFFFFFFFFFF000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000FFFFFFFFFFFF000000000000000000000000),
    .INIT_67(256'hFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFF000000000000),
    .INIT_68(256'hFFFFFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFF),
    .INIT_69(256'h0000FFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFF),
    .INIT_6A(256'hFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFFFFFF00000000000000000000),
    .INIT_6B(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF),
    .INIT_6C(256'h000000000000000000000000FFFFFFFFFFFF0000000000000000000000000000),
    .INIT_6D(256'hFFFFFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000),
    .INIT_6E(256'hFFFF0000000000000000000000000000FFFFFFFFFFFF0000000000000000FFFF),
    .INIT_6F(256'h0000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000FFFFFFFF),
    .INIT_70(256'hFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000),
    .INIT_71(256'hFFFFFFFFFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000),
    .INIT_72(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_73(256'hFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_74(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFF),
    .INIT_75(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_76(256'h000000000000000000000000FFFFFFFFFFFF0000000000000000000000000000),
    .INIT_77(256'hFFFFFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000),
    .INIT_78(256'hFFFF0000000000000000000000000000FFFFFFFFFFFF0000000000000000FFFF),
    .INIT_79(256'h0000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000FFFFFFFF),
    .INIT_7A(256'hFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000),
    .INIT_7B(256'hFFFFFFFFFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000),
    .INIT_7C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_7D(256'hFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_7E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFF),
    .INIT_7F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_20480x16_sub_016384_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_Naddra[12]_Naddr_o_al_n16 ),
    .dia({open_n507,open_n508,open_n509,open_n510,open_n511,open_n512,open_n513,open_n514,dia[7:0]}),
    .wea(wea),
    .doa({open_n536,open_n537,open_n538,open_n539,open_n540,open_n541,open_n542,open_n543,inst_doa_i4_007,inst_doa_i4_006,inst_doa_i4_005,inst_doa_i4_004,inst_doa_i4_003,inst_doa_i4_002,inst_doa_i4_001,inst_doa_i4_000}));
  // address_offset=16384;data_offset=8;depth=4096;width=8;num_section=1;width_per_section=8;section_size=16;working_depth=4096;working_width=8;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h000000000000FFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFF00000000),
    .INIT_02(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'h000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFF),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFF0FFFFFFFFFFFFFF7F7F7F7F7F3F3F1F1F0F030000),
    .INIT_09(256'h0F0300000000030F1F1F3F3F7F7F7F7F7FFFFFFFFFFFFFFFF0FFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000030F1F1F3F3F7F7F7F7F3F3F1F1F),
    .INIT_0B(256'h7FFFFFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFF7F7F7F7F3F3F3F1F0F07030000000003070F1F3F3F3F7F7F7F),
    .INIT_0D(256'h7F7F7F7F7FFFFFFFFFFFFFF0F0FFFFFFFFFFFF7F7F7F7F7F3F3F1F1F0F030000),
    .INIT_0E(256'h0F0300000000030F1F1F3F3F7F7F7F7F3F3F1F1F0F0300000000030F1F1F3F3F),
    .INIT_0F(256'hFFFFFFFFFFFFFEFEFEFCFCF8F8F0E0C00000030F1F1F3F3F7F7F7F7F3F3F1F1F),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFCFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFF7F7F3F1F0F0300000000030F1F3F7F7FFFFFC0E0F0F8F8FCFCFEFEFEFFFF),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h000000000000000000008080C0C0F0FCFCF0C0C0808000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h00000000000000000000000000008080C0C0F0FCFCF0C0C08080000000000000),
    .INIT_17(256'h0000000000008080C0C0F0FCFCF0C0C080800000000000000000000000000000),
    .INIT_18(256'h00000000FCF0C0C0808000000000000000008080C0C0F0F00000000000000000),
    .INIT_19(256'h808000000000000000008080C0C0F0FCFCF0C0C0808000000000000000000000),
    .INIT_1A(256'h00008080C0C0F0FCFCF0C0C0808000000000000000008080C0C0F0FCFCF0C0C0),
    .INIT_1B(256'hFCF0C0C0808000000000000000008080C0C0F0FC000000000000000000000000),
    .INIT_1C(256'h3C3C3C3C3C3C3F3F00000000000000003F3F30303030303030303F3F00000000),
    .INIT_1D(256'h00000000000000003F3F3F3F3F3F3F3F3F3F3F3F00000000000000003F3F3C3C),
    .INIT_1E(256'h3F3F3F3F3F3F3F3F3F3F3F3F00000000000000003F3F3F3F3F3F3F3F3F3F3F3F),
    .INIT_1F(256'h3F3F3F3F00000000000000003F3F3F3F3F3F3F3F3F3F3F3F0000000000000000),
    .INIT_20(256'h00000000FFFF0000000000000000FFFF00000000000000003F3F3F3F3F3F3F3F),
    .INIT_21(256'hF0F0F0F0F0F0FFFF0000000000000000FFFFC0C0C0C0C0C0C0C0FFFF00000000),
    .INIT_22(256'h0000000000000000FFFFFCFCFCFCFCFCFCFCFFFF0000000000000000FFFFF0F0),
    .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_24(256'hFFFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
    .INIT_25(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF),
    .INIT_26(256'hC0C0C0C0C0C0FFFF0000000000000000FFFF0000000000000000FFFF00000000),
    .INIT_27(256'h0000000000000000FFFFF0F0F0F0F0F0F0F0FFFF0000000000000000FFFFC0C0),
    .INIT_28(256'hFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000FFFFFCFCFCFCFCFCFCFCFFFF),
    .INIT_29(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h00000000000000003F3F3F3F0000000000000000000000000000000000000000),
    .INIT_31(256'h3F3F3F3F00000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h000000003F3F3F3F3F3F00000000000000000000000000000000000000000000),
    .INIT_33(256'h3F3F00000000000000000000000000003F3F3F3F3F3F00003F3F3F3F00000000),
    .INIT_34(256'h00000000000000003F3F3F3F3F3F00003F3F3F3F00000000000000003F3F3F3F),
    .INIT_35(256'h00000000000000003F3F3F3F0000000000000000000000000000000000000000),
    .INIT_36(256'h3F3F3F3F00000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h000000003F3F3F3F3F3F00000000000000000000000000000000000000000000),
    .INIT_38(256'h3F3F00000000000000000000000000003F3F3F3F3F3F00003F3F3F3F00000000),
    .INIT_39(256'h00000000000000003F3F3F3F3F3F00003F3F3F3F00000000000000003F3F3F3F),
    .INIT_3A(256'h00000000000000003F3F3F3F00003F3F3F3F0000000000000000000000000000),
    .INIT_3B(256'h3F3F3F3F00003F3F3F3F000000000000000000000000000000003F3F3F3F0000),
    .INIT_3C(256'h3F3F00003F3F3F3F3F3F00000000000000003F3F3F3F00000000000000000000),
    .INIT_3D(256'h3F3F00000000000000003F3F3F3F00003F3F3F3F3F3F00003F3F3F3F00003F3F),
    .INIT_3E(256'h00003F3F3F3F00003F3F3F3F3F3F00003F3F3F3F00003F3F3F3F00003F3F3F3F),
    .INIT_3F(256'h00000000000000003F3F3F3F00003F3F3F3F0000000000000000000000000000),
    .INIT_40(256'h3F3F3F3F00003F3F3F3F000000000000000000000000000000003F3F3F3F0000),
    .INIT_41(256'h3F3F00003F3F3F3F3F3F00000000000000003F3F3F3F00000000000000000000),
    .INIT_42(256'h3F3F00000000000000003F3F3F3F00003F3F3F3F3F3F00003F3F3F3F00003F3F),
    .INIT_43(256'h00003F3F3F3F00003F3F3F3F3F3F00003F3F3F3F00003F3F3F3F00003F3F3F3F),
    .INIT_44(256'h00000000000000003F3F3F3F0000000000000000000000000000000000000000),
    .INIT_45(256'h3F3F3F3F00000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h000000003F3F3F3F3F3F00000000000000000000000000000000000000000000),
    .INIT_47(256'h3F3F00000000000000000000000000003F3F3F3F3F3F00003F3F3F3F00000000),
    .INIT_48(256'h00000000000000003F3F3F3F3F3F00003F3F3F3F00000000000000003F3F3F3F),
    .INIT_49(256'h00000000000000003F3F3F3F0000000000000000000000000000000000000000),
    .INIT_4A(256'h3F3F3F3F00000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h000000003F3F3F3F3F3F00000000000000000000000000000000000000000000),
    .INIT_4C(256'h3F3F00000000000000000000000000003F3F3F3F3F3F00003F3F3F3F00000000),
    .INIT_4D(256'h00000000000000003F3F3F3F3F3F00003F3F3F3F00000000000000003F3F3F3F),
    .INIT_4E(256'h00000000000000003F3F3F3F00003F3F3F3F0000000000000000000000000000),
    .INIT_4F(256'h3F3F3F3F00003F3F3F3F000000000000000000000000000000003F3F3F3F0000),
    .INIT_50(256'h3F3F00003F3F3F3F3F3F00000000000000003F3F3F3F00000000000000000000),
    .INIT_51(256'h3F3F00000000000000003F3F3F3F00003F3F3F3F3F3F00003F3F3F3F00003F3F),
    .INIT_52(256'h00003F3F3F3F00003F3F3F3F3F3F00003F3F3F3F00003F3F3F3F00003F3F3F3F),
    .INIT_53(256'h00000000000000003F3F3F3F00003F3F3F3F0000000000000000000000000000),
    .INIT_54(256'h3F3F3F3F00003F3F3F3F000000000000000000000000000000003F3F3F3F0000),
    .INIT_55(256'h3F3F00003F3F3F3F3F3F00000000000000003F3F3F3F00000000000000000000),
    .INIT_56(256'h3F3F00000000000000003F3F3F3F00003F3F3F3F3F3F00003F3F3F3F00003F3F),
    .INIT_57(256'h00003F3F3F3F00003F3F3F3F3F3F00003F3F3F3F00003F3F3F3F00003F3F3F3F),
    .INIT_58(256'h000000000000FFFFFFFFFFFF0000000000000000000000000000000000000000),
    .INIT_59(256'hFFFFFFFF00000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000FFFFFFFFFFFFFFFF0000000000000000000000000000000000000000FFFF),
    .INIT_5B(256'hFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000),
    .INIT_5C(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF),
    .INIT_5D(256'h000000000000FFFFFFFFFFFF0000000000000000000000000000000000000000),
    .INIT_5E(256'hFFFFFFFF00000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000FFFFFFFFFFFFFFFF0000000000000000000000000000000000000000FFFF),
    .INIT_60(256'hFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000),
    .INIT_61(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF),
    .INIT_62(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000),
    .INIT_63(256'hFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000FFFFFFFFFFFF0000),
    .INIT_64(256'hFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF0000000000000000FFFF),
    .INIT_65(256'hFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_66(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_67(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000),
    .INIT_68(256'hFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000FFFFFFFFFFFF0000),
    .INIT_69(256'hFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF0000000000000000FFFF),
    .INIT_6A(256'hFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6C(256'h000000000000FFFFFFFFFFFF0000000000000000000000000000000000000000),
    .INIT_6D(256'hFFFFFFFF00000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000FFFFFFFFFFFFFFFF0000000000000000000000000000000000000000FFFF),
    .INIT_6F(256'hFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000),
    .INIT_70(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF),
    .INIT_71(256'h000000000000FFFFFFFFFFFF0000000000000000000000000000000000000000),
    .INIT_72(256'hFFFFFFFF00000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000FFFFFFFFFFFFFFFF0000000000000000000000000000000000000000FFFF),
    .INIT_74(256'hFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000),
    .INIT_75(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF),
    .INIT_76(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000),
    .INIT_77(256'hFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000FFFFFFFFFFFF0000),
    .INIT_78(256'hFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF0000000000000000FFFF),
    .INIT_79(256'hFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_7A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_7B(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000),
    .INIT_7C(256'hFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000FFFFFFFFFFFF0000),
    .INIT_7D(256'hFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFF0000000000000000FFFF),
    .INIT_7E(256'hFFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_7F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_20480x16_sub_016384_008 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_Naddra[12]_Naddr_o_al_n16 ),
    .dia({open_n564,open_n565,open_n566,open_n567,open_n568,open_n569,open_n570,open_n571,dia[15:8]}),
    .wea(wea),
    .doa({open_n593,open_n594,open_n595,open_n596,open_n597,open_n598,open_n599,open_n600,inst_doa_i4_015,inst_doa_i4_014,inst_doa_i4_013,inst_doa_i4_012,inst_doa_i4_011,inst_doa_i4_010,inst_doa_i4_009,inst_doa_i4_008}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b0/B1_0 ),
    .i1(inst_doa_i4_000),
    .sel(addra_piped[2]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b1/B1_0 ),
    .i1(inst_doa_i4_001),
    .sel(addra_piped[2]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_0  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i1_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_1  (
    .i0(inst_doa_i2_010),
    .i1(inst_doa_i3_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b10/B0_0 ),
    .i1(\inst_doa_mux_b10/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b10/B1_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b10/B1_0 ),
    .i1(inst_doa_i4_010),
    .sel(addra_piped[2]),
    .o(doa[10]));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_0  (
    .i0(inst_doa_i0_011),
    .i1(inst_doa_i1_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_1  (
    .i0(inst_doa_i2_011),
    .i1(inst_doa_i3_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b11/B0_0 ),
    .i1(\inst_doa_mux_b11/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b11/B1_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b11/B1_0 ),
    .i1(inst_doa_i4_011),
    .sel(addra_piped[2]),
    .o(doa[11]));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_0  (
    .i0(inst_doa_i0_012),
    .i1(inst_doa_i1_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_0 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_1  (
    .i0(inst_doa_i2_012),
    .i1(inst_doa_i3_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_1 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b12/B0_0 ),
    .i1(\inst_doa_mux_b12/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b12/B1_0 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b12/B1_0 ),
    .i1(inst_doa_i4_012),
    .sel(addra_piped[2]),
    .o(doa[12]));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_0  (
    .i0(inst_doa_i0_013),
    .i1(inst_doa_i1_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_0 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_1  (
    .i0(inst_doa_i2_013),
    .i1(inst_doa_i3_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_1 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b13/B0_0 ),
    .i1(\inst_doa_mux_b13/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b13/B1_0 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b13/B1_0 ),
    .i1(inst_doa_i4_013),
    .sel(addra_piped[2]),
    .o(doa[13]));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_0  (
    .i0(inst_doa_i0_014),
    .i1(inst_doa_i1_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_0 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_1  (
    .i0(inst_doa_i2_014),
    .i1(inst_doa_i3_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_1 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b14/B0_0 ),
    .i1(\inst_doa_mux_b14/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b14/B1_0 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b14/B1_0 ),
    .i1(inst_doa_i4_014),
    .sel(addra_piped[2]),
    .o(doa[14]));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_0  (
    .i0(inst_doa_i0_015),
    .i1(inst_doa_i1_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_0 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_1  (
    .i0(inst_doa_i2_015),
    .i1(inst_doa_i3_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_1 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b15/B0_0 ),
    .i1(\inst_doa_mux_b15/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b15/B1_0 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b15/B1_0 ),
    .i1(inst_doa_i4_015),
    .sel(addra_piped[2]),
    .o(doa[15]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b2/B1_0 ),
    .i1(inst_doa_i4_002),
    .sel(addra_piped[2]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b3/B1_0 ),
    .i1(inst_doa_i4_003),
    .sel(addra_piped[2]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b4/B1_0 ),
    .i1(inst_doa_i4_004),
    .sel(addra_piped[2]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b5/B1_0 ),
    .i1(inst_doa_i4_005),
    .sel(addra_piped[2]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b6/B1_0 ),
    .i1(inst_doa_i4_006),
    .sel(addra_piped[2]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b7/B1_0 ),
    .i1(inst_doa_i4_007),
    .sel(addra_piped[2]),
    .o(doa[7]));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_0  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i1_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_1  (
    .i0(inst_doa_i2_008),
    .i1(inst_doa_i3_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b8/B0_0 ),
    .i1(\inst_doa_mux_b8/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b8/B1_0 ),
    .i1(inst_doa_i4_008),
    .sel(addra_piped[2]),
    .o(doa[8]));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_0  (
    .i0(inst_doa_i0_009),
    .i1(inst_doa_i1_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_1  (
    .i0(inst_doa_i2_009),
    .i1(inst_doa_i3_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b9/B0_0 ),
    .i1(\inst_doa_mux_b9/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b9/B1_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b9/B1_0 ),
    .i1(inst_doa_i4_009),
    .sel(addra_piped[2]),
    .o(doa[9]));
  not wea_inv (wea_neg, wea);

endmodule 

module AL_DFF_X
  (
  ar,
  as,
  clk,
  d,
  en,
  sr,
  ss,
  q
  );

  input ar;
  input as;
  input clk;
  input d;
  input en;
  input sr;
  input ss;
  output q;

  wire enout;
  wire srout;
  wire ssout;

  AL_MUX u_en (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset (
    .i0(ssout),
    .i1(1'b0),
    .sel(sr),
    .o(srout));
  AL_DFF u_seq (
    .clk(clk),
    .d(srout),
    .reset(ar),
    .set(as),
    .q(q));
  AL_MUX u_set (
    .i0(enout),
    .i1(1'b1),
    .sel(ss),
    .o(ssout));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  // synthesis translate_off
  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end
  // synthesis translate_on

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule


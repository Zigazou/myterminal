module font (
	input wire clk,
	input wire [14:0] font_address,
	output reg [15:0] char_row_bitmap
);

reg [29:0] fifo = 30'd0;
always @(posedge clk) fifo <= { font_address, fifo[29:15] };

always @(posedge clk)
    case (fifo[14:0])
		15'h0000: char_row_bitmap <= 16'b0000000000000000;
		15'h0001: char_row_bitmap <= 16'b0000000000000000;
		15'h0002: char_row_bitmap <= 16'b0000111111000000;
		15'h0003: char_row_bitmap <= 16'b0001111111100000;
		15'h0004: char_row_bitmap <= 16'b0011100001110000;
		15'h0005: char_row_bitmap <= 16'b0011000000110000;
		15'h0006: char_row_bitmap <= 16'b0011000000000000;
		15'h0007: char_row_bitmap <= 16'b0011100000000000;
		15'h0008: char_row_bitmap <= 16'b0001110000000000;
		15'h0009: char_row_bitmap <= 16'b0000111000000000;
		15'h000a: char_row_bitmap <= 16'b0000011100000000;
		15'h000b: char_row_bitmap <= 16'b0000001100000000;
		15'h000c: char_row_bitmap <= 16'b0000000000000000;
		15'h000d: char_row_bitmap <= 16'b0000000000000000;
		15'h000e: char_row_bitmap <= 16'b0000001100000000;
		15'h000f: char_row_bitmap <= 16'b0000001100000000;
		15'h0010: char_row_bitmap <= 16'b0000000000000000;
		15'h0011: char_row_bitmap <= 16'b0000000000000000;
		15'h0012: char_row_bitmap <= 16'b0000000000000000;
		15'h0013: char_row_bitmap <= 16'b0000000000000000;
		15'h0014: char_row_bitmap <= 16'b0000000000000000;
		15'h0015: char_row_bitmap <= 16'b0000000000000000;
		15'h0016: char_row_bitmap <= 16'b0000001100000000;
		15'h0017: char_row_bitmap <= 16'b0000011110000000;
		15'h0018: char_row_bitmap <= 16'b0000111111000000;
		15'h0019: char_row_bitmap <= 16'b0000110011000000;
		15'h001a: char_row_bitmap <= 16'b0000000000000000;
		15'h001b: char_row_bitmap <= 16'b0000000000000000;
		15'h001c: char_row_bitmap <= 16'b0000111111000000;
		15'h001d: char_row_bitmap <= 16'b0001111111100000;
		15'h001e: char_row_bitmap <= 16'b0011100001110000;
		15'h001f: char_row_bitmap <= 16'b0011000000110000;
		15'h0020: char_row_bitmap <= 16'b0011111111110000;
		15'h0021: char_row_bitmap <= 16'b0011111111110000;
		15'h0022: char_row_bitmap <= 16'b0011000000110000;
		15'h0023: char_row_bitmap <= 16'b0011000000110000;
		15'h0024: char_row_bitmap <= 16'b0000000000000000;
		15'h0025: char_row_bitmap <= 16'b0000000000000000;
		15'h0026: char_row_bitmap <= 16'b0000000000000000;
		15'h0027: char_row_bitmap <= 16'b0000000000000000;
		15'h0028: char_row_bitmap <= 16'b0000000000000000;
		15'h0029: char_row_bitmap <= 16'b0000000011000000;
		15'h002a: char_row_bitmap <= 16'b0000000111000000;
		15'h002b: char_row_bitmap <= 16'b0000001110000000;
		15'h002c: char_row_bitmap <= 16'b0000001100000000;
		15'h002d: char_row_bitmap <= 16'b0000000000000000;
		15'h002e: char_row_bitmap <= 16'b0000111111110000;
		15'h002f: char_row_bitmap <= 16'b0000111111110000;
		15'h0030: char_row_bitmap <= 16'b0000110000000000;
		15'h0031: char_row_bitmap <= 16'b0000110000000000;
		15'h0032: char_row_bitmap <= 16'b0000111100000000;
		15'h0033: char_row_bitmap <= 16'b0000111100000000;
		15'h0034: char_row_bitmap <= 16'b0000110000000000;
		15'h0035: char_row_bitmap <= 16'b0000110000000000;
		15'h0036: char_row_bitmap <= 16'b0000111111110000;
		15'h0037: char_row_bitmap <= 16'b0000111111110000;
		15'h0038: char_row_bitmap <= 16'b0000000000000000;
		15'h0039: char_row_bitmap <= 16'b0000000000000000;
		15'h003a: char_row_bitmap <= 16'b0000000000000000;
		15'h003b: char_row_bitmap <= 16'b0000000000000000;
		15'h003c: char_row_bitmap <= 16'b0000000000000000;
		15'h003d: char_row_bitmap <= 16'b0000000000000000;
		15'h003e: char_row_bitmap <= 16'b0000000011000000;
		15'h003f: char_row_bitmap <= 16'b0000000111100000;
		15'h0040: char_row_bitmap <= 16'b0000001111110000;
		15'h0041: char_row_bitmap <= 16'b0000001100110000;
		15'h0042: char_row_bitmap <= 16'b0000001100000000;
		15'h0043: char_row_bitmap <= 16'b0000001100000000;
		15'h0044: char_row_bitmap <= 16'b0000111111000000;
		15'h0045: char_row_bitmap <= 16'b0000111111000000;
		15'h0046: char_row_bitmap <= 16'b0000001100000000;
		15'h0047: char_row_bitmap <= 16'b0000011100000000;
		15'h0048: char_row_bitmap <= 16'b0000111000110000;
		15'h0049: char_row_bitmap <= 16'b0000110000110000;
		15'h004a: char_row_bitmap <= 16'b0000111111110000;
		15'h004b: char_row_bitmap <= 16'b0000111111110000;
		15'h004c: char_row_bitmap <= 16'b0000000000000000;
		15'h004d: char_row_bitmap <= 16'b0000000000000000;
		15'h004e: char_row_bitmap <= 16'b0000000000000000;
		15'h004f: char_row_bitmap <= 16'b0000000000000000;
		15'h0050: char_row_bitmap <= 16'b0000000000000000;
		15'h0051: char_row_bitmap <= 16'b0000001100000000;
		15'h0052: char_row_bitmap <= 16'b0000011110000000;
		15'h0053: char_row_bitmap <= 16'b0000111111000000;
		15'h0054: char_row_bitmap <= 16'b0000110011000000;
		15'h0055: char_row_bitmap <= 16'b0000000000000000;
		15'h0056: char_row_bitmap <= 16'b0000111100110000;
		15'h0057: char_row_bitmap <= 16'b0001111110110000;
		15'h0058: char_row_bitmap <= 16'b0011100111110000;
		15'h0059: char_row_bitmap <= 16'b0011000011110000;
		15'h005a: char_row_bitmap <= 16'b0011000001110000;
		15'h005b: char_row_bitmap <= 16'b0011000001110000;
		15'h005c: char_row_bitmap <= 16'b0011000011110000;
		15'h005d: char_row_bitmap <= 16'b0011100111110000;
		15'h005e: char_row_bitmap <= 16'b0001111110110000;
		15'h005f: char_row_bitmap <= 16'b0000111100110000;
		15'h0060: char_row_bitmap <= 16'b0000000000000000;
		15'h0061: char_row_bitmap <= 16'b0000000000000000;
		15'h0062: char_row_bitmap <= 16'b0000000000000000;
		15'h0063: char_row_bitmap <= 16'b0000000000000000;
		15'h0064: char_row_bitmap <= 16'b0000000000000000;
		15'h0065: char_row_bitmap <= 16'b0000000000000000;
		15'h0066: char_row_bitmap <= 16'b0000111111000000;
		15'h0067: char_row_bitmap <= 16'b0001111111100000;
		15'h0068: char_row_bitmap <= 16'b0011100001110000;
		15'h0069: char_row_bitmap <= 16'b0011000000110000;
		15'h006a: char_row_bitmap <= 16'b0011000000000000;
		15'h006b: char_row_bitmap <= 16'b0011000000000000;
		15'h006c: char_row_bitmap <= 16'b0011000000000000;
		15'h006d: char_row_bitmap <= 16'b0011000000000000;
		15'h006e: char_row_bitmap <= 16'b0011000000000000;
		15'h006f: char_row_bitmap <= 16'b0011000000000000;
		15'h0070: char_row_bitmap <= 16'b0011000000110000;
		15'h0071: char_row_bitmap <= 16'b0011100001110000;
		15'h0072: char_row_bitmap <= 16'b0001111111100000;
		15'h0073: char_row_bitmap <= 16'b0000111111000000;
		15'h0074: char_row_bitmap <= 16'b0000001100000000;
		15'h0075: char_row_bitmap <= 16'b0000011100000000;
		15'h0076: char_row_bitmap <= 16'b0000111000000000;
		15'h0077: char_row_bitmap <= 16'b0000110000000000;
		15'h0078: char_row_bitmap <= 16'b0000000000000000;
		15'h0079: char_row_bitmap <= 16'b0000000000000000;
		15'h007a: char_row_bitmap <= 16'b0000011001100000;
		15'h007b: char_row_bitmap <= 16'b0000011001100000;
		15'h007c: char_row_bitmap <= 16'b0000000000000000;
		15'h007d: char_row_bitmap <= 16'b0000000000000000;
		15'h007e: char_row_bitmap <= 16'b0000111111110000;
		15'h007f: char_row_bitmap <= 16'b0000111111110000;
		15'h0080: char_row_bitmap <= 16'b0000110000000000;
		15'h0081: char_row_bitmap <= 16'b0000110000000000;
		15'h0082: char_row_bitmap <= 16'b0000111100000000;
		15'h0083: char_row_bitmap <= 16'b0000111100000000;
		15'h0084: char_row_bitmap <= 16'b0000110000000000;
		15'h0085: char_row_bitmap <= 16'b0000110000000000;
		15'h0086: char_row_bitmap <= 16'b0000111111110000;
		15'h0087: char_row_bitmap <= 16'b0000111111110000;
		15'h0088: char_row_bitmap <= 16'b0000000000000000;
		15'h0089: char_row_bitmap <= 16'b0000000000000000;
		15'h008a: char_row_bitmap <= 16'b0000000000000000;
		15'h008b: char_row_bitmap <= 16'b0000000000000000;
		15'h008c: char_row_bitmap <= 16'b0000000000000000;
		15'h008d: char_row_bitmap <= 16'b0000000000000000;
		15'h008e: char_row_bitmap <= 16'b0000110000000000;
		15'h008f: char_row_bitmap <= 16'b0000111000000000;
		15'h0090: char_row_bitmap <= 16'b0000011111000000;
		15'h0091: char_row_bitmap <= 16'b0000001111000000;
		15'h0092: char_row_bitmap <= 16'b0000000000000000;
		15'h0093: char_row_bitmap <= 16'b0000000000000000;
		15'h0094: char_row_bitmap <= 16'b0000111111000000;
		15'h0095: char_row_bitmap <= 16'b0001111111100000;
		15'h0096: char_row_bitmap <= 16'b0011100001110000;
		15'h0097: char_row_bitmap <= 16'b0011000000110000;
		15'h0098: char_row_bitmap <= 16'b0011111111110000;
		15'h0099: char_row_bitmap <= 16'b0011111111110000;
		15'h009a: char_row_bitmap <= 16'b0011000000110000;
		15'h009b: char_row_bitmap <= 16'b0011000000110000;
		15'h009c: char_row_bitmap <= 16'b0000000000000000;
		15'h009d: char_row_bitmap <= 16'b0000000000000000;
		15'h009e: char_row_bitmap <= 16'b0000000000000000;
		15'h009f: char_row_bitmap <= 16'b0000000000000000;
		15'h00a0: char_row_bitmap <= 16'b0000000000000000;
		15'h00a1: char_row_bitmap <= 16'b0000000000000000;
		15'h00a2: char_row_bitmap <= 16'b0000110000000000;
		15'h00a3: char_row_bitmap <= 16'b0000111000000000;
		15'h00a4: char_row_bitmap <= 16'b0000011111000000;
		15'h00a5: char_row_bitmap <= 16'b0000001111000000;
		15'h00a6: char_row_bitmap <= 16'b0000000000000000;
		15'h00a7: char_row_bitmap <= 16'b0000000000000000;
		15'h00a8: char_row_bitmap <= 16'b0011000000110000;
		15'h00a9: char_row_bitmap <= 16'b0011000000110000;
		15'h00aa: char_row_bitmap <= 16'b0011000000110000;
		15'h00ab: char_row_bitmap <= 16'b0011000001110000;
		15'h00ac: char_row_bitmap <= 16'b0011000011110000;
		15'h00ad: char_row_bitmap <= 16'b0011100111110000;
		15'h00ae: char_row_bitmap <= 16'b0001111110110000;
		15'h00af: char_row_bitmap <= 16'b0000111100110000;
		15'h00b0: char_row_bitmap <= 16'b0000000000000000;
		15'h00b1: char_row_bitmap <= 16'b0000000000000000;
		15'h00b2: char_row_bitmap <= 16'b0000000000000000;
		15'h00b3: char_row_bitmap <= 16'b0000000000000000;
		15'h00b4: char_row_bitmap <= 16'b0000000000000000;
		15'h00b5: char_row_bitmap <= 16'b0000001100000000;
		15'h00b6: char_row_bitmap <= 16'b0000001110000000;
		15'h00b7: char_row_bitmap <= 16'b0000000111000000;
		15'h00b8: char_row_bitmap <= 16'b0000000011000000;
		15'h00b9: char_row_bitmap <= 16'b0000000000000000;
		15'h00ba: char_row_bitmap <= 16'b0000111111110000;
		15'h00bb: char_row_bitmap <= 16'b0000111111110000;
		15'h00bc: char_row_bitmap <= 16'b0000110000000000;
		15'h00bd: char_row_bitmap <= 16'b0000110000000000;
		15'h00be: char_row_bitmap <= 16'b0000111100000000;
		15'h00bf: char_row_bitmap <= 16'b0000111100000000;
		15'h00c0: char_row_bitmap <= 16'b0000110000000000;
		15'h00c1: char_row_bitmap <= 16'b0000110000000000;
		15'h00c2: char_row_bitmap <= 16'b0000111111110000;
		15'h00c3: char_row_bitmap <= 16'b0000111111110000;
		15'h00c4: char_row_bitmap <= 16'b0000000000000000;
		15'h00c5: char_row_bitmap <= 16'b0000000000000000;
		15'h00c6: char_row_bitmap <= 16'b0000000000000000;
		15'h00c7: char_row_bitmap <= 16'b0000000000000000;
		15'h00c8: char_row_bitmap <= 16'b0000000000000000;
		15'h00c9: char_row_bitmap <= 16'b0000000000000000;
		15'h00ca: char_row_bitmap <= 16'b0000111111110000;
		15'h00cb: char_row_bitmap <= 16'b0001111111110000;
		15'h00cc: char_row_bitmap <= 16'b0011101100000000;
		15'h00cd: char_row_bitmap <= 16'b0011001100000000;
		15'h00ce: char_row_bitmap <= 16'b0011001100000000;
		15'h00cf: char_row_bitmap <= 16'b0011001100000000;
		15'h00d0: char_row_bitmap <= 16'b0011001111000000;
		15'h00d1: char_row_bitmap <= 16'b0011001111000000;
		15'h00d2: char_row_bitmap <= 16'b0011001100000000;
		15'h00d3: char_row_bitmap <= 16'b0011001100000000;
		15'h00d4: char_row_bitmap <= 16'b0011001100000000;
		15'h00d5: char_row_bitmap <= 16'b0011101100000000;
		15'h00d6: char_row_bitmap <= 16'b0001111111110000;
		15'h00d7: char_row_bitmap <= 16'b0000111111110000;
		15'h00d8: char_row_bitmap <= 16'b0000000000000000;
		15'h00d9: char_row_bitmap <= 16'b0000000000000000;
		15'h00da: char_row_bitmap <= 16'b0000000000000000;
		15'h00db: char_row_bitmap <= 16'b0000000000000000;
		15'h00dc: char_row_bitmap <= 16'b0000000000000000;
		15'h00dd: char_row_bitmap <= 16'b0000000011000000;
		15'h00de: char_row_bitmap <= 16'b0000000111100000;
		15'h00df: char_row_bitmap <= 16'b0000001111110000;
		15'h00e0: char_row_bitmap <= 16'b0000001100110000;
		15'h00e1: char_row_bitmap <= 16'b0000000000000000;
		15'h00e2: char_row_bitmap <= 16'b0000111111110000;
		15'h00e3: char_row_bitmap <= 16'b0000111111110000;
		15'h00e4: char_row_bitmap <= 16'b0000110000000000;
		15'h00e5: char_row_bitmap <= 16'b0000110000000000;
		15'h00e6: char_row_bitmap <= 16'b0000111100000000;
		15'h00e7: char_row_bitmap <= 16'b0000111100000000;
		15'h00e8: char_row_bitmap <= 16'b0000110000000000;
		15'h00e9: char_row_bitmap <= 16'b0000110000000000;
		15'h00ea: char_row_bitmap <= 16'b0000111111110000;
		15'h00eb: char_row_bitmap <= 16'b0000111111110000;
		15'h00ec: char_row_bitmap <= 16'b0000000000000000;
		15'h00ed: char_row_bitmap <= 16'b0000000000000000;
		15'h00ee: char_row_bitmap <= 16'b0000000000000000;
		15'h00ef: char_row_bitmap <= 16'b0000000000000000;
		15'h00f0: char_row_bitmap <= 16'b0000000000000000;
		15'h00f1: char_row_bitmap <= 16'b0000000000000000;
		15'h00f2: char_row_bitmap <= 16'b0000001111000000;
		15'h00f3: char_row_bitmap <= 16'b0000011111100000;
		15'h00f4: char_row_bitmap <= 16'b0000111001110000;
		15'h00f5: char_row_bitmap <= 16'b0000110000110000;
		15'h00f6: char_row_bitmap <= 16'b0011111110000000;
		15'h00f7: char_row_bitmap <= 16'b0011111110000000;
		15'h00f8: char_row_bitmap <= 16'b0000110000000000;
		15'h00f9: char_row_bitmap <= 16'b0000110000000000;
		15'h00fa: char_row_bitmap <= 16'b0011111110000000;
		15'h00fb: char_row_bitmap <= 16'b0011111110000000;
		15'h00fc: char_row_bitmap <= 16'b0000110000110000;
		15'h00fd: char_row_bitmap <= 16'b0000111001110000;
		15'h00fe: char_row_bitmap <= 16'b0000011111100000;
		15'h00ff: char_row_bitmap <= 16'b0000001111000000;
		15'h0100: char_row_bitmap <= 16'b0000000000000000;
		15'h0101: char_row_bitmap <= 16'b0000000000000000;
		15'h0102: char_row_bitmap <= 16'b0000000000000000;
		15'h0103: char_row_bitmap <= 16'b0000000000000000;
		15'h0104: char_row_bitmap <= 16'b0000000000000000;
		15'h0105: char_row_bitmap <= 16'b0000000000000000;
		15'h0106: char_row_bitmap <= 16'b0000001100000000;
		15'h0107: char_row_bitmap <= 16'b0000011110000000;
		15'h0108: char_row_bitmap <= 16'b0000111111000000;
		15'h0109: char_row_bitmap <= 16'b0000110011000000;
		15'h010a: char_row_bitmap <= 16'b0000000000000000;
		15'h010b: char_row_bitmap <= 16'b0000000000000000;
		15'h010c: char_row_bitmap <= 16'b0000111100000000;
		15'h010d: char_row_bitmap <= 16'b0000111100000000;
		15'h010e: char_row_bitmap <= 16'b0000001100000000;
		15'h010f: char_row_bitmap <= 16'b0000001100000000;
		15'h0110: char_row_bitmap <= 16'b0000001100000000;
		15'h0111: char_row_bitmap <= 16'b0000001100000000;
		15'h0112: char_row_bitmap <= 16'b0000111111000000;
		15'h0113: char_row_bitmap <= 16'b0000111111000000;
		15'h0114: char_row_bitmap <= 16'b0000000000000000;
		15'h0115: char_row_bitmap <= 16'b0000000000000000;
		15'h0116: char_row_bitmap <= 16'b0000000000000000;
		15'h0117: char_row_bitmap <= 16'b0000000000000000;
		15'h0118: char_row_bitmap <= 16'b0000000000000000;
		15'h0119: char_row_bitmap <= 16'b0000000000000000;
		15'h011a: char_row_bitmap <= 16'b0000011111100000;
		15'h011b: char_row_bitmap <= 16'b0001111111111000;
		15'h011c: char_row_bitmap <= 16'b0011110000111100;
		15'h011d: char_row_bitmap <= 16'b0011000000001100;
		15'h011e: char_row_bitmap <= 16'b0111001111001110;
		15'h011f: char_row_bitmap <= 16'b0110011111000110;
		15'h0120: char_row_bitmap <= 16'b0110011000000110;
		15'h0121: char_row_bitmap <= 16'b0110011000000110;
		15'h0122: char_row_bitmap <= 16'b0110011000000110;
		15'h0123: char_row_bitmap <= 16'b0110011000000110;
		15'h0124: char_row_bitmap <= 16'b0110011111000110;
		15'h0125: char_row_bitmap <= 16'b0111001111001110;
		15'h0126: char_row_bitmap <= 16'b0011000000001100;
		15'h0127: char_row_bitmap <= 16'b0011110000111100;
		15'h0128: char_row_bitmap <= 16'b0001111111111000;
		15'h0129: char_row_bitmap <= 16'b0000011111100000;
		15'h012a: char_row_bitmap <= 16'b0000000000000000;
		15'h012b: char_row_bitmap <= 16'b0000000000000000;
		15'h012c: char_row_bitmap <= 16'b0000000000000000;
		15'h012d: char_row_bitmap <= 16'b0000000000000000;
		15'h012e: char_row_bitmap <= 16'b0000011111100000;
		15'h012f: char_row_bitmap <= 16'b0001111111111000;
		15'h0130: char_row_bitmap <= 16'b0011110000111100;
		15'h0131: char_row_bitmap <= 16'b0011000000001100;
		15'h0132: char_row_bitmap <= 16'b0111011111001110;
		15'h0133: char_row_bitmap <= 16'b0110011111100110;
		15'h0134: char_row_bitmap <= 16'b0110011001100110;
		15'h0135: char_row_bitmap <= 16'b0110011111100110;
		15'h0136: char_row_bitmap <= 16'b0110011111000110;
		15'h0137: char_row_bitmap <= 16'b0110011011000110;
		15'h0138: char_row_bitmap <= 16'b0110011001100110;
		15'h0139: char_row_bitmap <= 16'b0111011001101110;
		15'h013a: char_row_bitmap <= 16'b0011000000001100;
		15'h013b: char_row_bitmap <= 16'b0011110000111100;
		15'h013c: char_row_bitmap <= 16'b0001111111111000;
		15'h013d: char_row_bitmap <= 16'b0000011111100000;
		15'h013e: char_row_bitmap <= 16'b0000000000000000;
		15'h013f: char_row_bitmap <= 16'b0000000000000000;
		15'h0140: char_row_bitmap <= 16'b0000000000000000;
		15'h0141: char_row_bitmap <= 16'b0000000000000000;
		15'h0142: char_row_bitmap <= 16'b0000001110000000;
		15'h0143: char_row_bitmap <= 16'b0000011111000000;
		15'h0144: char_row_bitmap <= 16'b0000111011100000;
		15'h0145: char_row_bitmap <= 16'b0000110001100000;
		15'h0146: char_row_bitmap <= 16'b0000111011100000;
		15'h0147: char_row_bitmap <= 16'b0000011111000000;
		15'h0148: char_row_bitmap <= 16'b0000001110000000;
		15'h0149: char_row_bitmap <= 16'b0000000000000000;
		15'h014a: char_row_bitmap <= 16'b0000000000000000;
		15'h014b: char_row_bitmap <= 16'b0000000000000000;
		15'h014c: char_row_bitmap <= 16'b0000000000000000;
		15'h014d: char_row_bitmap <= 16'b0000000000000000;
		15'h014e: char_row_bitmap <= 16'b0000000000000000;
		15'h014f: char_row_bitmap <= 16'b0000000000000000;
		15'h0150: char_row_bitmap <= 16'b0000000000000000;
		15'h0151: char_row_bitmap <= 16'b0000000000000000;
		15'h0152: char_row_bitmap <= 16'b0000000000000000;
		15'h0153: char_row_bitmap <= 16'b0000000000000000;
		15'h0154: char_row_bitmap <= 16'b0000000000000000;
		15'h0155: char_row_bitmap <= 16'b0000000000000000;
		15'h0156: char_row_bitmap <= 16'b0000001100000000;
		15'h0157: char_row_bitmap <= 16'b0000001100000000;
		15'h0158: char_row_bitmap <= 16'b0000001100000000;
		15'h0159: char_row_bitmap <= 16'b0000001100000000;
		15'h015a: char_row_bitmap <= 16'b0011111111110000;
		15'h015b: char_row_bitmap <= 16'b0011111111110000;
		15'h015c: char_row_bitmap <= 16'b0000001100000000;
		15'h015d: char_row_bitmap <= 16'b0000001100000000;
		15'h015e: char_row_bitmap <= 16'b0000001100000000;
		15'h015f: char_row_bitmap <= 16'b0000001100000000;
		15'h0160: char_row_bitmap <= 16'b0000000000000000;
		15'h0161: char_row_bitmap <= 16'b0000000000000000;
		15'h0162: char_row_bitmap <= 16'b0011111111110000;
		15'h0163: char_row_bitmap <= 16'b0011111111110000;
		15'h0164: char_row_bitmap <= 16'b0000000000000000;
		15'h0165: char_row_bitmap <= 16'b0000000000000000;
		15'h0166: char_row_bitmap <= 16'b0000000000000000;
		15'h0167: char_row_bitmap <= 16'b0000000000000000;
		15'h0168: char_row_bitmap <= 16'b0000000000000000;
		15'h0169: char_row_bitmap <= 16'b0000000011000000;
		15'h016a: char_row_bitmap <= 16'b0000000111000000;
		15'h016b: char_row_bitmap <= 16'b0000001110000000;
		15'h016c: char_row_bitmap <= 16'b0000001100000000;
		15'h016d: char_row_bitmap <= 16'b0000000000000000;
		15'h016e: char_row_bitmap <= 16'b0000111111000000;
		15'h016f: char_row_bitmap <= 16'b0001111111100000;
		15'h0170: char_row_bitmap <= 16'b0011100001110000;
		15'h0171: char_row_bitmap <= 16'b0011000000110000;
		15'h0172: char_row_bitmap <= 16'b0011111111110000;
		15'h0173: char_row_bitmap <= 16'b0011111111110000;
		15'h0174: char_row_bitmap <= 16'b0011000000000000;
		15'h0175: char_row_bitmap <= 16'b0011100000000000;
		15'h0176: char_row_bitmap <= 16'b0001111111100000;
		15'h0177: char_row_bitmap <= 16'b0000111111100000;
		15'h0178: char_row_bitmap <= 16'b0000000000000000;
		15'h0179: char_row_bitmap <= 16'b0000000000000000;
		15'h017a: char_row_bitmap <= 16'b0000000000000000;
		15'h017b: char_row_bitmap <= 16'b0000000000000000;
		15'h017c: char_row_bitmap <= 16'b0000000000000000;
		15'h017d: char_row_bitmap <= 16'b0000000000000000;
		15'h017e: char_row_bitmap <= 16'b0000110011000000;
		15'h017f: char_row_bitmap <= 16'b0000110011000000;
		15'h0180: char_row_bitmap <= 16'b0000000000000000;
		15'h0181: char_row_bitmap <= 16'b0000000000000000;
		15'h0182: char_row_bitmap <= 16'b0000111111000000;
		15'h0183: char_row_bitmap <= 16'b0001111111100000;
		15'h0184: char_row_bitmap <= 16'b0011100001110000;
		15'h0185: char_row_bitmap <= 16'b0011000000110000;
		15'h0186: char_row_bitmap <= 16'b0011111111110000;
		15'h0187: char_row_bitmap <= 16'b0011111111110000;
		15'h0188: char_row_bitmap <= 16'b0011000000000000;
		15'h0189: char_row_bitmap <= 16'b0011100000000000;
		15'h018a: char_row_bitmap <= 16'b0001111111100000;
		15'h018b: char_row_bitmap <= 16'b0000111111100000;
		15'h018c: char_row_bitmap <= 16'b0000000000000000;
		15'h018d: char_row_bitmap <= 16'b0000000000000000;
		15'h018e: char_row_bitmap <= 16'b0000000000000000;
		15'h018f: char_row_bitmap <= 16'b0000000000000000;
		15'h0190: char_row_bitmap <= 16'b0000000000000000;
		15'h0191: char_row_bitmap <= 16'b0000000000000000;
		15'h0192: char_row_bitmap <= 16'b0000110011000000;
		15'h0193: char_row_bitmap <= 16'b0000110011000000;
		15'h0194: char_row_bitmap <= 16'b0000000000000000;
		15'h0195: char_row_bitmap <= 16'b0000000000000000;
		15'h0196: char_row_bitmap <= 16'b0000111100000000;
		15'h0197: char_row_bitmap <= 16'b0000111100000000;
		15'h0198: char_row_bitmap <= 16'b0000001100000000;
		15'h0199: char_row_bitmap <= 16'b0000001100000000;
		15'h019a: char_row_bitmap <= 16'b0000001100000000;
		15'h019b: char_row_bitmap <= 16'b0000001100000000;
		15'h019c: char_row_bitmap <= 16'b0000001100000000;
		15'h019d: char_row_bitmap <= 16'b0000001100000000;
		15'h019e: char_row_bitmap <= 16'b0000111111000000;
		15'h019f: char_row_bitmap <= 16'b0000111111000000;
		15'h01a0: char_row_bitmap <= 16'b0000000000000000;
		15'h01a1: char_row_bitmap <= 16'b0000000000000000;
		15'h01a2: char_row_bitmap <= 16'b0000000000000000;
		15'h01a3: char_row_bitmap <= 16'b0000000000000000;
		15'h01a4: char_row_bitmap <= 16'b0000000000000000;
		15'h01a5: char_row_bitmap <= 16'b0000000000000000;
		15'h01a6: char_row_bitmap <= 16'b0000000000000000;
		15'h01a7: char_row_bitmap <= 16'b0000000000000000;
		15'h01a8: char_row_bitmap <= 16'b0000000000000000;
		15'h01a9: char_row_bitmap <= 16'b0000000000000000;
		15'h01aa: char_row_bitmap <= 16'b0000111111000000;
		15'h01ab: char_row_bitmap <= 16'b0001111111000000;
		15'h01ac: char_row_bitmap <= 16'b0011100000000000;
		15'h01ad: char_row_bitmap <= 16'b0011000000000000;
		15'h01ae: char_row_bitmap <= 16'b0011000000000000;
		15'h01af: char_row_bitmap <= 16'b0011000000000000;
		15'h01b0: char_row_bitmap <= 16'b0011000000000000;
		15'h01b1: char_row_bitmap <= 16'b0011100000000000;
		15'h01b2: char_row_bitmap <= 16'b0001111111000000;
		15'h01b3: char_row_bitmap <= 16'b0000111111000000;
		15'h01b4: char_row_bitmap <= 16'b0000001100000000;
		15'h01b5: char_row_bitmap <= 16'b0000011100000000;
		15'h01b6: char_row_bitmap <= 16'b0000111000000000;
		15'h01b7: char_row_bitmap <= 16'b0000110000000000;
		15'h01b8: char_row_bitmap <= 16'b0000000000000000;
		15'h01b9: char_row_bitmap <= 16'b0000000000000000;
		15'h01ba: char_row_bitmap <= 16'b0000001100000000;
		15'h01bb: char_row_bitmap <= 16'b0000011110000000;
		15'h01bc: char_row_bitmap <= 16'b0000111111000000;
		15'h01bd: char_row_bitmap <= 16'b0000110011000000;
		15'h01be: char_row_bitmap <= 16'b0000000000000000;
		15'h01bf: char_row_bitmap <= 16'b0000000000000000;
		15'h01c0: char_row_bitmap <= 16'b0011000000110000;
		15'h01c1: char_row_bitmap <= 16'b0011000000110000;
		15'h01c2: char_row_bitmap <= 16'b0011000000110000;
		15'h01c3: char_row_bitmap <= 16'b0011000001110000;
		15'h01c4: char_row_bitmap <= 16'b0011000011110000;
		15'h01c5: char_row_bitmap <= 16'b0011100111110000;
		15'h01c6: char_row_bitmap <= 16'b0001111110110000;
		15'h01c7: char_row_bitmap <= 16'b0000111100110000;
		15'h01c8: char_row_bitmap <= 16'b0000000000000000;
		15'h01c9: char_row_bitmap <= 16'b0000000000000000;
		15'h01ca: char_row_bitmap <= 16'b0000000000000000;
		15'h01cb: char_row_bitmap <= 16'b0000000000000000;
		15'h01cc: char_row_bitmap <= 16'b0000000000000000;
		15'h01cd: char_row_bitmap <= 16'b0000110000000000;
		15'h01ce: char_row_bitmap <= 16'b0000111000000000;
		15'h01cf: char_row_bitmap <= 16'b0000011100000000;
		15'h01d0: char_row_bitmap <= 16'b0000001100000000;
		15'h01d1: char_row_bitmap <= 16'b0000000000000000;
		15'h01d2: char_row_bitmap <= 16'b0000111100110000;
		15'h01d3: char_row_bitmap <= 16'b0001111110110000;
		15'h01d4: char_row_bitmap <= 16'b0011100111110000;
		15'h01d5: char_row_bitmap <= 16'b0011000011110000;
		15'h01d6: char_row_bitmap <= 16'b0011000001110000;
		15'h01d7: char_row_bitmap <= 16'b0011000001110000;
		15'h01d8: char_row_bitmap <= 16'b0011000011110000;
		15'h01d9: char_row_bitmap <= 16'b0011100111110000;
		15'h01da: char_row_bitmap <= 16'b0001111110110000;
		15'h01db: char_row_bitmap <= 16'b0000111100110000;
		15'h01dc: char_row_bitmap <= 16'b0000000000000000;
		15'h01dd: char_row_bitmap <= 16'b0000000000000000;
		15'h01de: char_row_bitmap <= 16'b0000000000000000;
		15'h01df: char_row_bitmap <= 16'b0000000000000000;
		15'h01e0: char_row_bitmap <= 16'b0000000000000000;
		15'h01e1: char_row_bitmap <= 16'b0000000000000000;
		15'h01e2: char_row_bitmap <= 16'b0000000000000000;
		15'h01e3: char_row_bitmap <= 16'b0000000000000000;
		15'h01e4: char_row_bitmap <= 16'b0000001100000000;
		15'h01e5: char_row_bitmap <= 16'b0000001100000000;
		15'h01e6: char_row_bitmap <= 16'b0000000000000000;
		15'h01e7: char_row_bitmap <= 16'b0000000000000000;
		15'h01e8: char_row_bitmap <= 16'b0011111111110000;
		15'h01e9: char_row_bitmap <= 16'b0011111111110000;
		15'h01ea: char_row_bitmap <= 16'b0000000000000000;
		15'h01eb: char_row_bitmap <= 16'b0000000000000000;
		15'h01ec: char_row_bitmap <= 16'b0000001100000000;
		15'h01ed: char_row_bitmap <= 16'b0000001100000000;
		15'h01ee: char_row_bitmap <= 16'b0000000000000000;
		15'h01ef: char_row_bitmap <= 16'b0000000000000000;
		15'h01f0: char_row_bitmap <= 16'b0000000000000000;
		15'h01f1: char_row_bitmap <= 16'b0000000000000000;
		15'h01f2: char_row_bitmap <= 16'b0000000000000000;
		15'h01f3: char_row_bitmap <= 16'b0000000000000000;
		15'h01f4: char_row_bitmap <= 16'b0000000000000000;
		15'h01f5: char_row_bitmap <= 16'b0000110000000000;
		15'h01f6: char_row_bitmap <= 16'b0000111000000000;
		15'h01f7: char_row_bitmap <= 16'b0000011100000000;
		15'h01f8: char_row_bitmap <= 16'b0000001100000000;
		15'h01f9: char_row_bitmap <= 16'b0000000000000000;
		15'h01fa: char_row_bitmap <= 16'b0000111111000000;
		15'h01fb: char_row_bitmap <= 16'b0001111111100000;
		15'h01fc: char_row_bitmap <= 16'b0011100001110000;
		15'h01fd: char_row_bitmap <= 16'b0011000000110000;
		15'h01fe: char_row_bitmap <= 16'b0011111111110000;
		15'h01ff: char_row_bitmap <= 16'b0011111111110000;
		15'h0200: char_row_bitmap <= 16'b0011000000000000;
		15'h0201: char_row_bitmap <= 16'b0011100000000000;
		15'h0202: char_row_bitmap <= 16'b0001111111100000;
		15'h0203: char_row_bitmap <= 16'b0000111111100000;
		15'h0204: char_row_bitmap <= 16'b0000000000000000;
		15'h0205: char_row_bitmap <= 16'b0000000000000000;
		15'h0206: char_row_bitmap <= 16'b0000000000000000;
		15'h0207: char_row_bitmap <= 16'b0000000000000000;
		15'h0208: char_row_bitmap <= 16'b0000000000000000;
		15'h0209: char_row_bitmap <= 16'b0000000000000000;
		15'h020a: char_row_bitmap <= 16'b0000000000000000;
		15'h020b: char_row_bitmap <= 16'b0000000000000000;
		15'h020c: char_row_bitmap <= 16'b0000000000000000;
		15'h020d: char_row_bitmap <= 16'b0000000000000000;
		15'h020e: char_row_bitmap <= 16'b0000111111110000;
		15'h020f: char_row_bitmap <= 16'b0001111111111000;
		15'h0210: char_row_bitmap <= 16'b0011101110011100;
		15'h0211: char_row_bitmap <= 16'b0011001100001100;
		15'h0212: char_row_bitmap <= 16'b0011001111111100;
		15'h0213: char_row_bitmap <= 16'b0011001111111100;
		15'h0214: char_row_bitmap <= 16'b0011001100000000;
		15'h0215: char_row_bitmap <= 16'b0011101100000000;
		15'h0216: char_row_bitmap <= 16'b0001111111111000;
		15'h0217: char_row_bitmap <= 16'b0000111111111000;
		15'h0218: char_row_bitmap <= 16'b0000000000000000;
		15'h0219: char_row_bitmap <= 16'b0000000000000000;
		15'h021a: char_row_bitmap <= 16'b0000000000000000;
		15'h021b: char_row_bitmap <= 16'b0000000000000000;
		15'h021c: char_row_bitmap <= 16'b0000000000000000;
		15'h021d: char_row_bitmap <= 16'b0000001100000000;
		15'h021e: char_row_bitmap <= 16'b0000011110000000;
		15'h021f: char_row_bitmap <= 16'b0000111111000000;
		15'h0220: char_row_bitmap <= 16'b0000110011000000;
		15'h0221: char_row_bitmap <= 16'b0000000000000000;
		15'h0222: char_row_bitmap <= 16'b0000111111000000;
		15'h0223: char_row_bitmap <= 16'b0001111111100000;
		15'h0224: char_row_bitmap <= 16'b0011100001110000;
		15'h0225: char_row_bitmap <= 16'b0011000000110000;
		15'h0226: char_row_bitmap <= 16'b0011111111110000;
		15'h0227: char_row_bitmap <= 16'b0011111111110000;
		15'h0228: char_row_bitmap <= 16'b0011000000000000;
		15'h0229: char_row_bitmap <= 16'b0011100000000000;
		15'h022a: char_row_bitmap <= 16'b0001111111100000;
		15'h022b: char_row_bitmap <= 16'b0000111111100000;
		15'h022c: char_row_bitmap <= 16'b0000000000000000;
		15'h022d: char_row_bitmap <= 16'b0000000000000000;
		15'h022e: char_row_bitmap <= 16'b0000000000000000;
		15'h022f: char_row_bitmap <= 16'b0000000000000000;
		15'h0230: char_row_bitmap <= 16'b0000000000000000;
		15'h0231: char_row_bitmap <= 16'b0000000000000000;
		15'h0232: char_row_bitmap <= 16'b0011000000000000;
		15'h0233: char_row_bitmap <= 16'b0111000000000000;
		15'h0234: char_row_bitmap <= 16'b1111000000000000;
		15'h0235: char_row_bitmap <= 16'b1111000000000000;
		15'h0236: char_row_bitmap <= 16'b0011000000000000;
		15'h0237: char_row_bitmap <= 16'b0011000000000000;
		15'h0238: char_row_bitmap <= 16'b0011000000110000;
		15'h0239: char_row_bitmap <= 16'b0011000001110000;
		15'h023a: char_row_bitmap <= 16'b0011000011110000;
		15'h023b: char_row_bitmap <= 16'b0011000111110000;
		15'h023c: char_row_bitmap <= 16'b0000001110110000;
		15'h023d: char_row_bitmap <= 16'b0000011100110000;
		15'h023e: char_row_bitmap <= 16'b0000011111111100;
		15'h023f: char_row_bitmap <= 16'b0000011111111100;
		15'h0240: char_row_bitmap <= 16'b0000000000110000;
		15'h0241: char_row_bitmap <= 16'b0000000000110000;
		15'h0242: char_row_bitmap <= 16'b0000000000000000;
		15'h0243: char_row_bitmap <= 16'b0000000000000000;
		15'h0244: char_row_bitmap <= 16'b0000000000000000;
		15'h0245: char_row_bitmap <= 16'b0000000000000000;
		15'h0246: char_row_bitmap <= 16'b0011000000000000;
		15'h0247: char_row_bitmap <= 16'b0111000000000000;
		15'h0248: char_row_bitmap <= 16'b1111000000000000;
		15'h0249: char_row_bitmap <= 16'b1111000000000000;
		15'h024a: char_row_bitmap <= 16'b0011000000000000;
		15'h024b: char_row_bitmap <= 16'b0011000000000000;
		15'h024c: char_row_bitmap <= 16'b0011000011110000;
		15'h024d: char_row_bitmap <= 16'b0011000111111000;
		15'h024e: char_row_bitmap <= 16'b0011001110011100;
		15'h024f: char_row_bitmap <= 16'b0011001100011100;
		15'h0250: char_row_bitmap <= 16'b0000000000111000;
		15'h0251: char_row_bitmap <= 16'b0000000001110000;
		15'h0252: char_row_bitmap <= 16'b0000000011100000;
		15'h0253: char_row_bitmap <= 16'b0000000111000000;
		15'h0254: char_row_bitmap <= 16'b0000001111111100;
		15'h0255: char_row_bitmap <= 16'b0000001111111100;
		15'h0256: char_row_bitmap <= 16'b0000000000000000;
		15'h0257: char_row_bitmap <= 16'b0000000000000000;
		15'h0258: char_row_bitmap <= 16'b0000000000000000;
		15'h0259: char_row_bitmap <= 16'b0000000000000000;
		15'h025a: char_row_bitmap <= 16'b1111000000000000;
		15'h025b: char_row_bitmap <= 16'b1111100000000000;
		15'h025c: char_row_bitmap <= 16'b0001110000000000;
		15'h025d: char_row_bitmap <= 16'b0001110000000000;
		15'h025e: char_row_bitmap <= 16'b0011100000000000;
		15'h025f: char_row_bitmap <= 16'b0011100000000000;
		15'h0260: char_row_bitmap <= 16'b0001110000110000;
		15'h0261: char_row_bitmap <= 16'b0001110001110000;
		15'h0262: char_row_bitmap <= 16'b1111100011110000;
		15'h0263: char_row_bitmap <= 16'b1111000111110000;
		15'h0264: char_row_bitmap <= 16'b0000001110110000;
		15'h0265: char_row_bitmap <= 16'b0000011100110000;
		15'h0266: char_row_bitmap <= 16'b0000011111111100;
		15'h0267: char_row_bitmap <= 16'b0000011111111100;
		15'h0268: char_row_bitmap <= 16'b0000000000110000;
		15'h0269: char_row_bitmap <= 16'b0000000000110000;
		15'h026a: char_row_bitmap <= 16'b0000000000000000;
		15'h026b: char_row_bitmap <= 16'b0000000000000000;
		15'h026c: char_row_bitmap <= 16'b0000000000000000;
		15'h026d: char_row_bitmap <= 16'b0000000000000000;
		15'h026e: char_row_bitmap <= 16'b0000001100000000;
		15'h026f: char_row_bitmap <= 16'b0000011110000000;
		15'h0270: char_row_bitmap <= 16'b0000111111000000;
		15'h0271: char_row_bitmap <= 16'b0000110011000000;
		15'h0272: char_row_bitmap <= 16'b0000000000000000;
		15'h0273: char_row_bitmap <= 16'b0000111111000000;
		15'h0274: char_row_bitmap <= 16'b0001111111100000;
		15'h0275: char_row_bitmap <= 16'b0011100001110000;
		15'h0276: char_row_bitmap <= 16'b0011000000110000;
		15'h0277: char_row_bitmap <= 16'b0011000000110000;
		15'h0278: char_row_bitmap <= 16'b0011000000110000;
		15'h0279: char_row_bitmap <= 16'b0011100001110000;
		15'h027a: char_row_bitmap <= 16'b0001111111100000;
		15'h027b: char_row_bitmap <= 16'b0000111111000000;
		15'h027c: char_row_bitmap <= 16'b0000000000000000;
		15'h027d: char_row_bitmap <= 16'b0000000000000000;
		15'h027e: char_row_bitmap <= 16'b0000000000000000;
		15'h027f: char_row_bitmap <= 16'b0000000000000000;
		15'h0280: char_row_bitmap <= 16'b0000000000000000;
		15'h0281: char_row_bitmap <= 16'b0000000000000000;
		15'h0282: char_row_bitmap <= 16'b0000000000000000;
		15'h0283: char_row_bitmap <= 16'b0000000000000000;
		15'h0284: char_row_bitmap <= 16'b0000000000000000;
		15'h0285: char_row_bitmap <= 16'b0000000000000000;
		15'h0286: char_row_bitmap <= 16'b0000000000000000;
		15'h0287: char_row_bitmap <= 16'b0000000000000000;
		15'h0288: char_row_bitmap <= 16'b0000000000000000;
		15'h0289: char_row_bitmap <= 16'b0000000000000000;
		15'h028a: char_row_bitmap <= 16'b0000000000000000;
		15'h028b: char_row_bitmap <= 16'b0000000000000000;
		15'h028c: char_row_bitmap <= 16'b0000000000000000;
		15'h028d: char_row_bitmap <= 16'b0000000000000000;
		15'h028e: char_row_bitmap <= 16'b0000000000000000;
		15'h028f: char_row_bitmap <= 16'b0000000000000000;
		15'h0290: char_row_bitmap <= 16'b0000000000000000;
		15'h0291: char_row_bitmap <= 16'b0000000000000000;
		15'h0292: char_row_bitmap <= 16'b0000000000000000;
		15'h0293: char_row_bitmap <= 16'b0000000000000000;
		15'h0294: char_row_bitmap <= 16'b0000000000000000;
		15'h0295: char_row_bitmap <= 16'b0000000000000000;
		15'h0296: char_row_bitmap <= 16'b0000001100000000;
		15'h0297: char_row_bitmap <= 16'b0000001100000000;
		15'h0298: char_row_bitmap <= 16'b0000001100000000;
		15'h0299: char_row_bitmap <= 16'b0000001100000000;
		15'h029a: char_row_bitmap <= 16'b0000001100000000;
		15'h029b: char_row_bitmap <= 16'b0000001100000000;
		15'h029c: char_row_bitmap <= 16'b0000001100000000;
		15'h029d: char_row_bitmap <= 16'b0000001100000000;
		15'h029e: char_row_bitmap <= 16'b0000001100000000;
		15'h029f: char_row_bitmap <= 16'b0000001100000000;
		15'h02a0: char_row_bitmap <= 16'b0000000000000000;
		15'h02a1: char_row_bitmap <= 16'b0000000000000000;
		15'h02a2: char_row_bitmap <= 16'b0000001100000000;
		15'h02a3: char_row_bitmap <= 16'b0000001100000000;
		15'h02a4: char_row_bitmap <= 16'b0000000000000000;
		15'h02a5: char_row_bitmap <= 16'b0000000000000000;
		15'h02a6: char_row_bitmap <= 16'b0000000000000000;
		15'h02a7: char_row_bitmap <= 16'b0000000000000000;
		15'h02a8: char_row_bitmap <= 16'b0000000000000000;
		15'h02a9: char_row_bitmap <= 16'b0000000000000000;
		15'h02aa: char_row_bitmap <= 16'b0000110011000000;
		15'h02ab: char_row_bitmap <= 16'b0000110011000000;
		15'h02ac: char_row_bitmap <= 16'b0000110011000000;
		15'h02ad: char_row_bitmap <= 16'b0000110011000000;
		15'h02ae: char_row_bitmap <= 16'b0000110011000000;
		15'h02af: char_row_bitmap <= 16'b0000110011000000;
		15'h02b0: char_row_bitmap <= 16'b0000000000000000;
		15'h02b1: char_row_bitmap <= 16'b0000000000000000;
		15'h02b2: char_row_bitmap <= 16'b0000000000000000;
		15'h02b3: char_row_bitmap <= 16'b0000000000000000;
		15'h02b4: char_row_bitmap <= 16'b0000000000000000;
		15'h02b5: char_row_bitmap <= 16'b0000000000000000;
		15'h02b6: char_row_bitmap <= 16'b0000000000000000;
		15'h02b7: char_row_bitmap <= 16'b0000000000000000;
		15'h02b8: char_row_bitmap <= 16'b0000000000000000;
		15'h02b9: char_row_bitmap <= 16'b0000000000000000;
		15'h02ba: char_row_bitmap <= 16'b0000000000000000;
		15'h02bb: char_row_bitmap <= 16'b0000000000000000;
		15'h02bc: char_row_bitmap <= 16'b0000000000000000;
		15'h02bd: char_row_bitmap <= 16'b0000000000000000;
		15'h02be: char_row_bitmap <= 16'b0000110011000000;
		15'h02bf: char_row_bitmap <= 16'b0000110011000000;
		15'h02c0: char_row_bitmap <= 16'b0000110011000000;
		15'h02c1: char_row_bitmap <= 16'b0000110011000000;
		15'h02c2: char_row_bitmap <= 16'b0011110011110000;
		15'h02c3: char_row_bitmap <= 16'b0011110011110000;
		15'h02c4: char_row_bitmap <= 16'b0000110011000000;
		15'h02c5: char_row_bitmap <= 16'b0000110011000000;
		15'h02c6: char_row_bitmap <= 16'b0011110011110000;
		15'h02c7: char_row_bitmap <= 16'b0011110011110000;
		15'h02c8: char_row_bitmap <= 16'b0000110011000000;
		15'h02c9: char_row_bitmap <= 16'b0000110011000000;
		15'h02ca: char_row_bitmap <= 16'b0000110011000000;
		15'h02cb: char_row_bitmap <= 16'b0000110011000000;
		15'h02cc: char_row_bitmap <= 16'b0000000000000000;
		15'h02cd: char_row_bitmap <= 16'b0000000000000000;
		15'h02ce: char_row_bitmap <= 16'b0000000000000000;
		15'h02cf: char_row_bitmap <= 16'b0000000000000000;
		15'h02d0: char_row_bitmap <= 16'b0000000000000000;
		15'h02d1: char_row_bitmap <= 16'b0000001100000000;
		15'h02d2: char_row_bitmap <= 16'b0000001100000000;
		15'h02d3: char_row_bitmap <= 16'b0000111111100000;
		15'h02d4: char_row_bitmap <= 16'b0001111111110000;
		15'h02d5: char_row_bitmap <= 16'b0011101100110000;
		15'h02d6: char_row_bitmap <= 16'b0011001100000000;
		15'h02d7: char_row_bitmap <= 16'b0011101100000000;
		15'h02d8: char_row_bitmap <= 16'b0001111111000000;
		15'h02d9: char_row_bitmap <= 16'b0000111111100000;
		15'h02da: char_row_bitmap <= 16'b0000001101110000;
		15'h02db: char_row_bitmap <= 16'b0000001100110000;
		15'h02dc: char_row_bitmap <= 16'b0011001100110000;
		15'h02dd: char_row_bitmap <= 16'b0011101101110000;
		15'h02de: char_row_bitmap <= 16'b0001111111100000;
		15'h02df: char_row_bitmap <= 16'b0000111111000000;
		15'h02e0: char_row_bitmap <= 16'b0000001100000000;
		15'h02e1: char_row_bitmap <= 16'b0000001100000000;
		15'h02e2: char_row_bitmap <= 16'b0000000000000000;
		15'h02e3: char_row_bitmap <= 16'b0000000000000000;
		15'h02e4: char_row_bitmap <= 16'b0000000000000000;
		15'h02e5: char_row_bitmap <= 16'b0000000000000000;
		15'h02e6: char_row_bitmap <= 16'b0001100000000000;
		15'h02e7: char_row_bitmap <= 16'b0011110000000000;
		15'h02e8: char_row_bitmap <= 16'b0011110000110000;
		15'h02e9: char_row_bitmap <= 16'b0001100001110000;
		15'h02ea: char_row_bitmap <= 16'b0000000011100000;
		15'h02eb: char_row_bitmap <= 16'b0000000111000000;
		15'h02ec: char_row_bitmap <= 16'b0000001110000000;
		15'h02ed: char_row_bitmap <= 16'b0000011100000000;
		15'h02ee: char_row_bitmap <= 16'b0000111000000000;
		15'h02ef: char_row_bitmap <= 16'b0001110000000000;
		15'h02f0: char_row_bitmap <= 16'b0011100001100000;
		15'h02f1: char_row_bitmap <= 16'b0011000011110000;
		15'h02f2: char_row_bitmap <= 16'b0000000011110000;
		15'h02f3: char_row_bitmap <= 16'b0000000001100000;
		15'h02f4: char_row_bitmap <= 16'b0000000000000000;
		15'h02f5: char_row_bitmap <= 16'b0000000000000000;
		15'h02f6: char_row_bitmap <= 16'b0000000000000000;
		15'h02f7: char_row_bitmap <= 16'b0000000000000000;
		15'h02f8: char_row_bitmap <= 16'b0000000000000000;
		15'h02f9: char_row_bitmap <= 16'b0000000000000000;
		15'h02fa: char_row_bitmap <= 16'b0000110000000000;
		15'h02fb: char_row_bitmap <= 16'b0001111000000000;
		15'h02fc: char_row_bitmap <= 16'b0011111100000000;
		15'h02fd: char_row_bitmap <= 16'b0011001100000000;
		15'h02fe: char_row_bitmap <= 16'b0011001100000000;
		15'h02ff: char_row_bitmap <= 16'b0011111100000000;
		15'h0300: char_row_bitmap <= 16'b0001111000000000;
		15'h0301: char_row_bitmap <= 16'b0001110000000000;
		15'h0302: char_row_bitmap <= 16'b0011111100110000;
		15'h0303: char_row_bitmap <= 16'b0011001111110000;
		15'h0304: char_row_bitmap <= 16'b0011000111100000;
		15'h0305: char_row_bitmap <= 16'b0011100111100000;
		15'h0306: char_row_bitmap <= 16'b0001111111110000;
		15'h0307: char_row_bitmap <= 16'b0000111100110000;
		15'h0308: char_row_bitmap <= 16'b0000000000000000;
		15'h0309: char_row_bitmap <= 16'b0000000000000000;
		15'h030a: char_row_bitmap <= 16'b0000000000000000;
		15'h030b: char_row_bitmap <= 16'b0000000000000000;
		15'h030c: char_row_bitmap <= 16'b0000000000000000;
		15'h030d: char_row_bitmap <= 16'b0000000000000000;
		15'h030e: char_row_bitmap <= 16'b0000001100000000;
		15'h030f: char_row_bitmap <= 16'b0000001100000000;
		15'h0310: char_row_bitmap <= 16'b0000001100000000;
		15'h0311: char_row_bitmap <= 16'b0000011100000000;
		15'h0312: char_row_bitmap <= 16'b0000111000000000;
		15'h0313: char_row_bitmap <= 16'b0000110000000000;
		15'h0314: char_row_bitmap <= 16'b0000000000000000;
		15'h0315: char_row_bitmap <= 16'b0000000000000000;
		15'h0316: char_row_bitmap <= 16'b0000000000000000;
		15'h0317: char_row_bitmap <= 16'b0000000000000000;
		15'h0318: char_row_bitmap <= 16'b0000000000000000;
		15'h0319: char_row_bitmap <= 16'b0000000000000000;
		15'h031a: char_row_bitmap <= 16'b0000000000000000;
		15'h031b: char_row_bitmap <= 16'b0000000000000000;
		15'h031c: char_row_bitmap <= 16'b0000000000000000;
		15'h031d: char_row_bitmap <= 16'b0000000000000000;
		15'h031e: char_row_bitmap <= 16'b0000000000000000;
		15'h031f: char_row_bitmap <= 16'b0000000000000000;
		15'h0320: char_row_bitmap <= 16'b0000000000000000;
		15'h0321: char_row_bitmap <= 16'b0000000000000000;
		15'h0322: char_row_bitmap <= 16'b0000000011000000;
		15'h0323: char_row_bitmap <= 16'b0000000111000000;
		15'h0324: char_row_bitmap <= 16'b0000001110000000;
		15'h0325: char_row_bitmap <= 16'b0000011100000000;
		15'h0326: char_row_bitmap <= 16'b0000111000000000;
		15'h0327: char_row_bitmap <= 16'b0000110000000000;
		15'h0328: char_row_bitmap <= 16'b0000110000000000;
		15'h0329: char_row_bitmap <= 16'b0000110000000000;
		15'h032a: char_row_bitmap <= 16'b0000110000000000;
		15'h032b: char_row_bitmap <= 16'b0000110000000000;
		15'h032c: char_row_bitmap <= 16'b0000111000000000;
		15'h032d: char_row_bitmap <= 16'b0000011100000000;
		15'h032e: char_row_bitmap <= 16'b0000001110000000;
		15'h032f: char_row_bitmap <= 16'b0000000111000000;
		15'h0330: char_row_bitmap <= 16'b0000000011000000;
		15'h0331: char_row_bitmap <= 16'b0000000000000000;
		15'h0332: char_row_bitmap <= 16'b0000000000000000;
		15'h0333: char_row_bitmap <= 16'b0000000000000000;
		15'h0334: char_row_bitmap <= 16'b0000000000000000;
		15'h0335: char_row_bitmap <= 16'b0000000000000000;
		15'h0336: char_row_bitmap <= 16'b0000110000000000;
		15'h0337: char_row_bitmap <= 16'b0000111000000000;
		15'h0338: char_row_bitmap <= 16'b0000011100000000;
		15'h0339: char_row_bitmap <= 16'b0000001110000000;
		15'h033a: char_row_bitmap <= 16'b0000000111000000;
		15'h033b: char_row_bitmap <= 16'b0000000011000000;
		15'h033c: char_row_bitmap <= 16'b0000000011000000;
		15'h033d: char_row_bitmap <= 16'b0000000011000000;
		15'h033e: char_row_bitmap <= 16'b0000000011000000;
		15'h033f: char_row_bitmap <= 16'b0000000011000000;
		15'h0340: char_row_bitmap <= 16'b0000000111000000;
		15'h0341: char_row_bitmap <= 16'b0000001110000000;
		15'h0342: char_row_bitmap <= 16'b0000011100000000;
		15'h0343: char_row_bitmap <= 16'b0000111000000000;
		15'h0344: char_row_bitmap <= 16'b0000110000000000;
		15'h0345: char_row_bitmap <= 16'b0000000000000000;
		15'h0346: char_row_bitmap <= 16'b0000000000000000;
		15'h0347: char_row_bitmap <= 16'b0000000000000000;
		15'h0348: char_row_bitmap <= 16'b0000000000000000;
		15'h0349: char_row_bitmap <= 16'b0000000000000000;
		15'h034a: char_row_bitmap <= 16'b0000000000000000;
		15'h034b: char_row_bitmap <= 16'b0000001100000000;
		15'h034c: char_row_bitmap <= 16'b0011001100110000;
		15'h034d: char_row_bitmap <= 16'b0011101101110000;
		15'h034e: char_row_bitmap <= 16'b0001111111100000;
		15'h034f: char_row_bitmap <= 16'b0000111111000000;
		15'h0350: char_row_bitmap <= 16'b0000011110000000;
		15'h0351: char_row_bitmap <= 16'b0000011110000000;
		15'h0352: char_row_bitmap <= 16'b0000111111000000;
		15'h0353: char_row_bitmap <= 16'b0001111111100000;
		15'h0354: char_row_bitmap <= 16'b0011101101110000;
		15'h0355: char_row_bitmap <= 16'b0011001100110000;
		15'h0356: char_row_bitmap <= 16'b0000001100000000;
		15'h0357: char_row_bitmap <= 16'b0000000000000000;
		15'h0358: char_row_bitmap <= 16'b0000000000000000;
		15'h0359: char_row_bitmap <= 16'b0000000000000000;
		15'h035a: char_row_bitmap <= 16'b0000000000000000;
		15'h035b: char_row_bitmap <= 16'b0000000000000000;
		15'h035c: char_row_bitmap <= 16'b0000000000000000;
		15'h035d: char_row_bitmap <= 16'b0000000000000000;
		15'h035e: char_row_bitmap <= 16'b0000000000000000;
		15'h035f: char_row_bitmap <= 16'b0000000000000000;
		15'h0360: char_row_bitmap <= 16'b0000001100000000;
		15'h0361: char_row_bitmap <= 16'b0000001100000000;
		15'h0362: char_row_bitmap <= 16'b0000001100000000;
		15'h0363: char_row_bitmap <= 16'b0000001100000000;
		15'h0364: char_row_bitmap <= 16'b0011111111110000;
		15'h0365: char_row_bitmap <= 16'b0011111111110000;
		15'h0366: char_row_bitmap <= 16'b0000001100000000;
		15'h0367: char_row_bitmap <= 16'b0000001100000000;
		15'h0368: char_row_bitmap <= 16'b0000001100000000;
		15'h0369: char_row_bitmap <= 16'b0000001100000000;
		15'h036a: char_row_bitmap <= 16'b0000000000000000;
		15'h036b: char_row_bitmap <= 16'b0000000000000000;
		15'h036c: char_row_bitmap <= 16'b0000000000000000;
		15'h036d: char_row_bitmap <= 16'b0000000000000000;
		15'h036e: char_row_bitmap <= 16'b0000000000000000;
		15'h036f: char_row_bitmap <= 16'b0000000000000000;
		15'h0370: char_row_bitmap <= 16'b0000000000000000;
		15'h0371: char_row_bitmap <= 16'b0000000000000000;
		15'h0372: char_row_bitmap <= 16'b0000000000000000;
		15'h0373: char_row_bitmap <= 16'b0000000000000000;
		15'h0374: char_row_bitmap <= 16'b0000000000000000;
		15'h0375: char_row_bitmap <= 16'b0000000000000000;
		15'h0376: char_row_bitmap <= 16'b0000000000000000;
		15'h0377: char_row_bitmap <= 16'b0000000000000000;
		15'h0378: char_row_bitmap <= 16'b0000000000000000;
		15'h0379: char_row_bitmap <= 16'b0000000000000000;
		15'h037a: char_row_bitmap <= 16'b0000000000000000;
		15'h037b: char_row_bitmap <= 16'b0000000000000000;
		15'h037c: char_row_bitmap <= 16'b0000110000000000;
		15'h037d: char_row_bitmap <= 16'b0000110000000000;
		15'h037e: char_row_bitmap <= 16'b0000110000000000;
		15'h037f: char_row_bitmap <= 16'b0001110000000000;
		15'h0380: char_row_bitmap <= 16'b0011100000000000;
		15'h0381: char_row_bitmap <= 16'b0011000000000000;
		15'h0382: char_row_bitmap <= 16'b0000000000000000;
		15'h0383: char_row_bitmap <= 16'b0000000000000000;
		15'h0384: char_row_bitmap <= 16'b0000000000000000;
		15'h0385: char_row_bitmap <= 16'b0000000000000000;
		15'h0386: char_row_bitmap <= 16'b0000000000000000;
		15'h0387: char_row_bitmap <= 16'b0000000000000000;
		15'h0388: char_row_bitmap <= 16'b0000000000000000;
		15'h0389: char_row_bitmap <= 16'b0000000000000000;
		15'h038a: char_row_bitmap <= 16'b0000000000000000;
		15'h038b: char_row_bitmap <= 16'b0000000000000000;
		15'h038c: char_row_bitmap <= 16'b0000000000000000;
		15'h038d: char_row_bitmap <= 16'b0000000000000000;
		15'h038e: char_row_bitmap <= 16'b0000111111110000;
		15'h038f: char_row_bitmap <= 16'b0000111111110000;
		15'h0390: char_row_bitmap <= 16'b0000000000000000;
		15'h0391: char_row_bitmap <= 16'b0000000000000000;
		15'h0392: char_row_bitmap <= 16'b0000000000000000;
		15'h0393: char_row_bitmap <= 16'b0000000000000000;
		15'h0394: char_row_bitmap <= 16'b0000000000000000;
		15'h0395: char_row_bitmap <= 16'b0000000000000000;
		15'h0396: char_row_bitmap <= 16'b0000000000000000;
		15'h0397: char_row_bitmap <= 16'b0000000000000000;
		15'h0398: char_row_bitmap <= 16'b0000000000000000;
		15'h0399: char_row_bitmap <= 16'b0000000000000000;
		15'h039a: char_row_bitmap <= 16'b0000000000000000;
		15'h039b: char_row_bitmap <= 16'b0000000000000000;
		15'h039c: char_row_bitmap <= 16'b0000000000000000;
		15'h039d: char_row_bitmap <= 16'b0000000000000000;
		15'h039e: char_row_bitmap <= 16'b0000000000000000;
		15'h039f: char_row_bitmap <= 16'b0000000000000000;
		15'h03a0: char_row_bitmap <= 16'b0000000000000000;
		15'h03a1: char_row_bitmap <= 16'b0000000000000000;
		15'h03a2: char_row_bitmap <= 16'b0000000000000000;
		15'h03a3: char_row_bitmap <= 16'b0000000000000000;
		15'h03a4: char_row_bitmap <= 16'b0000000000000000;
		15'h03a5: char_row_bitmap <= 16'b0000000000000000;
		15'h03a6: char_row_bitmap <= 16'b0000110000000000;
		15'h03a7: char_row_bitmap <= 16'b0000110000000000;
		15'h03a8: char_row_bitmap <= 16'b0000000000000000;
		15'h03a9: char_row_bitmap <= 16'b0000000000000000;
		15'h03aa: char_row_bitmap <= 16'b0000000000000000;
		15'h03ab: char_row_bitmap <= 16'b0000000000000000;
		15'h03ac: char_row_bitmap <= 16'b0000000000000011;
		15'h03ad: char_row_bitmap <= 16'b0000000000000111;
		15'h03ae: char_row_bitmap <= 16'b0000000000000110;
		15'h03af: char_row_bitmap <= 16'b0000000000001100;
		15'h03b0: char_row_bitmap <= 16'b0000000000011100;
		15'h03b1: char_row_bitmap <= 16'b0000000000111000;
		15'h03b2: char_row_bitmap <= 16'b0000000001110000;
		15'h03b3: char_row_bitmap <= 16'b0000000001100000;
		15'h03b4: char_row_bitmap <= 16'b0000000011100000;
		15'h03b5: char_row_bitmap <= 16'b0000000111000000;
		15'h03b6: char_row_bitmap <= 16'b0000001110000000;
		15'h03b7: char_row_bitmap <= 16'b0000011100000000;
		15'h03b8: char_row_bitmap <= 16'b0000011000000000;
		15'h03b9: char_row_bitmap <= 16'b0000111000000000;
		15'h03ba: char_row_bitmap <= 16'b0001110000000000;
		15'h03bb: char_row_bitmap <= 16'b0011100000000000;
		15'h03bc: char_row_bitmap <= 16'b0111000000000000;
		15'h03bd: char_row_bitmap <= 16'b0110000000000000;
		15'h03be: char_row_bitmap <= 16'b1110000000000000;
		15'h03bf: char_row_bitmap <= 16'b1100000000000000;
		15'h03c0: char_row_bitmap <= 16'b0000000000000000;
		15'h03c1: char_row_bitmap <= 16'b0000000000000000;
		15'h03c2: char_row_bitmap <= 16'b0000001100000000;
		15'h03c3: char_row_bitmap <= 16'b0000011110000000;
		15'h03c4: char_row_bitmap <= 16'b0000111111000000;
		15'h03c5: char_row_bitmap <= 16'b0001110011100000;
		15'h03c6: char_row_bitmap <= 16'b0011100001110000;
		15'h03c7: char_row_bitmap <= 16'b0011000000110000;
		15'h03c8: char_row_bitmap <= 16'b0011000000110000;
		15'h03c9: char_row_bitmap <= 16'b0011000000110000;
		15'h03ca: char_row_bitmap <= 16'b0011000000110000;
		15'h03cb: char_row_bitmap <= 16'b0011100001110000;
		15'h03cc: char_row_bitmap <= 16'b0001110011100000;
		15'h03cd: char_row_bitmap <= 16'b0000111111000000;
		15'h03ce: char_row_bitmap <= 16'b0000011110000000;
		15'h03cf: char_row_bitmap <= 16'b0000001100000000;
		15'h03d0: char_row_bitmap <= 16'b0000000000000000;
		15'h03d1: char_row_bitmap <= 16'b0000000000000000;
		15'h03d2: char_row_bitmap <= 16'b0000000000000000;
		15'h03d3: char_row_bitmap <= 16'b0000000000000000;
		15'h03d4: char_row_bitmap <= 16'b0000000000000000;
		15'h03d5: char_row_bitmap <= 16'b0000000000000000;
		15'h03d6: char_row_bitmap <= 16'b0000001100000000;
		15'h03d7: char_row_bitmap <= 16'b0000011100000000;
		15'h03d8: char_row_bitmap <= 16'b0000111100000000;
		15'h03d9: char_row_bitmap <= 16'b0001111100000000;
		15'h03da: char_row_bitmap <= 16'b0000001100000000;
		15'h03db: char_row_bitmap <= 16'b0000001100000000;
		15'h03dc: char_row_bitmap <= 16'b0000001100000000;
		15'h03dd: char_row_bitmap <= 16'b0000001100000000;
		15'h03de: char_row_bitmap <= 16'b0000001100000000;
		15'h03df: char_row_bitmap <= 16'b0000001100000000;
		15'h03e0: char_row_bitmap <= 16'b0000001100000000;
		15'h03e1: char_row_bitmap <= 16'b0000001100000000;
		15'h03e2: char_row_bitmap <= 16'b0000001100000000;
		15'h03e3: char_row_bitmap <= 16'b0000001100000000;
		15'h03e4: char_row_bitmap <= 16'b0000000000000000;
		15'h03e5: char_row_bitmap <= 16'b0000000000000000;
		15'h03e6: char_row_bitmap <= 16'b0000000000000000;
		15'h03e7: char_row_bitmap <= 16'b0000000000000000;
		15'h03e8: char_row_bitmap <= 16'b0000000000000000;
		15'h03e9: char_row_bitmap <= 16'b0000000000000000;
		15'h03ea: char_row_bitmap <= 16'b0000111111000000;
		15'h03eb: char_row_bitmap <= 16'b0001111111100000;
		15'h03ec: char_row_bitmap <= 16'b0011100001110000;
		15'h03ed: char_row_bitmap <= 16'b0011000000110000;
		15'h03ee: char_row_bitmap <= 16'b0000000000110000;
		15'h03ef: char_row_bitmap <= 16'b0000000001110000;
		15'h03f0: char_row_bitmap <= 16'b0000001111100000;
		15'h03f1: char_row_bitmap <= 16'b0000011111000000;
		15'h03f2: char_row_bitmap <= 16'b0000111000000000;
		15'h03f3: char_row_bitmap <= 16'b0001110000000000;
		15'h03f4: char_row_bitmap <= 16'b0011100000000000;
		15'h03f5: char_row_bitmap <= 16'b0011000000000000;
		15'h03f6: char_row_bitmap <= 16'b0011111111110000;
		15'h03f7: char_row_bitmap <= 16'b0011111111110000;
		15'h03f8: char_row_bitmap <= 16'b0000000000000000;
		15'h03f9: char_row_bitmap <= 16'b0000000000000000;
		15'h03fa: char_row_bitmap <= 16'b0000000000000000;
		15'h03fb: char_row_bitmap <= 16'b0000000000000000;
		15'h03fc: char_row_bitmap <= 16'b0000000000000000;
		15'h03fd: char_row_bitmap <= 16'b0000000000000000;
		15'h03fe: char_row_bitmap <= 16'b0011111111110000;
		15'h03ff: char_row_bitmap <= 16'b0011111111110000;
		15'h0400: char_row_bitmap <= 16'b0000000000110000;
		15'h0401: char_row_bitmap <= 16'b0000000001110000;
		15'h0402: char_row_bitmap <= 16'b0000000011100000;
		15'h0403: char_row_bitmap <= 16'b0000000111000000;
		15'h0404: char_row_bitmap <= 16'b0000001111000000;
		15'h0405: char_row_bitmap <= 16'b0000001111100000;
		15'h0406: char_row_bitmap <= 16'b0000000001110000;
		15'h0407: char_row_bitmap <= 16'b0000000000110000;
		15'h0408: char_row_bitmap <= 16'b0011000000110000;
		15'h0409: char_row_bitmap <= 16'b0011100001110000;
		15'h040a: char_row_bitmap <= 16'b0001111111100000;
		15'h040b: char_row_bitmap <= 16'b0000111111000000;
		15'h040c: char_row_bitmap <= 16'b0000000000000000;
		15'h040d: char_row_bitmap <= 16'b0000000000000000;
		15'h040e: char_row_bitmap <= 16'b0000000000000000;
		15'h040f: char_row_bitmap <= 16'b0000000000000000;
		15'h0410: char_row_bitmap <= 16'b0000000000000000;
		15'h0411: char_row_bitmap <= 16'b0000000000000000;
		15'h0412: char_row_bitmap <= 16'b0000000011000000;
		15'h0413: char_row_bitmap <= 16'b0000000111000000;
		15'h0414: char_row_bitmap <= 16'b0000001111000000;
		15'h0415: char_row_bitmap <= 16'b0000011111000000;
		15'h0416: char_row_bitmap <= 16'b0000111011000000;
		15'h0417: char_row_bitmap <= 16'b0001110011000000;
		15'h0418: char_row_bitmap <= 16'b0011100011000000;
		15'h0419: char_row_bitmap <= 16'b0011000011000000;
		15'h041a: char_row_bitmap <= 16'b0011111111110000;
		15'h041b: char_row_bitmap <= 16'b0011111111110000;
		15'h041c: char_row_bitmap <= 16'b0000000011000000;
		15'h041d: char_row_bitmap <= 16'b0000000011000000;
		15'h041e: char_row_bitmap <= 16'b0000000011000000;
		15'h041f: char_row_bitmap <= 16'b0000000011000000;
		15'h0420: char_row_bitmap <= 16'b0000000000000000;
		15'h0421: char_row_bitmap <= 16'b0000000000000000;
		15'h0422: char_row_bitmap <= 16'b0000000000000000;
		15'h0423: char_row_bitmap <= 16'b0000000000000000;
		15'h0424: char_row_bitmap <= 16'b0000000000000000;
		15'h0425: char_row_bitmap <= 16'b0000000000000000;
		15'h0426: char_row_bitmap <= 16'b0011111111110000;
		15'h0427: char_row_bitmap <= 16'b0011111111110000;
		15'h0428: char_row_bitmap <= 16'b0011000000000000;
		15'h0429: char_row_bitmap <= 16'b0011000000000000;
		15'h042a: char_row_bitmap <= 16'b0011111111000000;
		15'h042b: char_row_bitmap <= 16'b0011111111100000;
		15'h042c: char_row_bitmap <= 16'b0000000001110000;
		15'h042d: char_row_bitmap <= 16'b0000000000110000;
		15'h042e: char_row_bitmap <= 16'b0000000000110000;
		15'h042f: char_row_bitmap <= 16'b0000000000110000;
		15'h0430: char_row_bitmap <= 16'b0011000000110000;
		15'h0431: char_row_bitmap <= 16'b0011100001110000;
		15'h0432: char_row_bitmap <= 16'b0001111111100000;
		15'h0433: char_row_bitmap <= 16'b0000111111000000;
		15'h0434: char_row_bitmap <= 16'b0000000000000000;
		15'h0435: char_row_bitmap <= 16'b0000000000000000;
		15'h0436: char_row_bitmap <= 16'b0000000000000000;
		15'h0437: char_row_bitmap <= 16'b0000000000000000;
		15'h0438: char_row_bitmap <= 16'b0000000000000000;
		15'h0439: char_row_bitmap <= 16'b0000000000000000;
		15'h043a: char_row_bitmap <= 16'b0000001111000000;
		15'h043b: char_row_bitmap <= 16'b0000011111000000;
		15'h043c: char_row_bitmap <= 16'b0000111000000000;
		15'h043d: char_row_bitmap <= 16'b0001110000000000;
		15'h043e: char_row_bitmap <= 16'b0011100000000000;
		15'h043f: char_row_bitmap <= 16'b0011000000000000;
		15'h0440: char_row_bitmap <= 16'b0011011111000000;
		15'h0441: char_row_bitmap <= 16'b0011111111100000;
		15'h0442: char_row_bitmap <= 16'b0011100001110000;
		15'h0443: char_row_bitmap <= 16'b0011000000110000;
		15'h0444: char_row_bitmap <= 16'b0011000000110000;
		15'h0445: char_row_bitmap <= 16'b0011100001110000;
		15'h0446: char_row_bitmap <= 16'b0001111111100000;
		15'h0447: char_row_bitmap <= 16'b0000111111000000;
		15'h0448: char_row_bitmap <= 16'b0000000000000000;
		15'h0449: char_row_bitmap <= 16'b0000000000000000;
		15'h044a: char_row_bitmap <= 16'b0000000000000000;
		15'h044b: char_row_bitmap <= 16'b0000000000000000;
		15'h044c: char_row_bitmap <= 16'b0000000000000000;
		15'h044d: char_row_bitmap <= 16'b0000000000000000;
		15'h044e: char_row_bitmap <= 16'b0011111111110000;
		15'h044f: char_row_bitmap <= 16'b0011111111110000;
		15'h0450: char_row_bitmap <= 16'b0000000000110000;
		15'h0451: char_row_bitmap <= 16'b0000000001110000;
		15'h0452: char_row_bitmap <= 16'b0000000011100000;
		15'h0453: char_row_bitmap <= 16'b0000000111000000;
		15'h0454: char_row_bitmap <= 16'b0000001110000000;
		15'h0455: char_row_bitmap <= 16'b0000011100000000;
		15'h0456: char_row_bitmap <= 16'b0000111000000000;
		15'h0457: char_row_bitmap <= 16'b0000110000000000;
		15'h0458: char_row_bitmap <= 16'b0000110000000000;
		15'h0459: char_row_bitmap <= 16'b0000110000000000;
		15'h045a: char_row_bitmap <= 16'b0000110000000000;
		15'h045b: char_row_bitmap <= 16'b0000110000000000;
		15'h045c: char_row_bitmap <= 16'b0000000000000000;
		15'h045d: char_row_bitmap <= 16'b0000000000000000;
		15'h045e: char_row_bitmap <= 16'b0000000000000000;
		15'h045f: char_row_bitmap <= 16'b0000000000000000;
		15'h0460: char_row_bitmap <= 16'b0000000000000000;
		15'h0461: char_row_bitmap <= 16'b0000000000000000;
		15'h0462: char_row_bitmap <= 16'b0000111111000000;
		15'h0463: char_row_bitmap <= 16'b0001111111100000;
		15'h0464: char_row_bitmap <= 16'b0011100001110000;
		15'h0465: char_row_bitmap <= 16'b0011000000110000;
		15'h0466: char_row_bitmap <= 16'b0011000000110000;
		15'h0467: char_row_bitmap <= 16'b0011000001110000;
		15'h0468: char_row_bitmap <= 16'b0001111111100000;
		15'h0469: char_row_bitmap <= 16'b0001111111100000;
		15'h046a: char_row_bitmap <= 16'b0011100001110000;
		15'h046b: char_row_bitmap <= 16'b0011000000110000;
		15'h046c: char_row_bitmap <= 16'b0011000000110000;
		15'h046d: char_row_bitmap <= 16'b0011100001110000;
		15'h046e: char_row_bitmap <= 16'b0001111111100000;
		15'h046f: char_row_bitmap <= 16'b0000111111000000;
		15'h0470: char_row_bitmap <= 16'b0000000000000000;
		15'h0471: char_row_bitmap <= 16'b0000000000000000;
		15'h0472: char_row_bitmap <= 16'b0000000000000000;
		15'h0473: char_row_bitmap <= 16'b0000000000000000;
		15'h0474: char_row_bitmap <= 16'b0000000000000000;
		15'h0475: char_row_bitmap <= 16'b0000000000000000;
		15'h0476: char_row_bitmap <= 16'b0000111111000000;
		15'h0477: char_row_bitmap <= 16'b0001111111100000;
		15'h0478: char_row_bitmap <= 16'b0011100001110000;
		15'h0479: char_row_bitmap <= 16'b0011000000110000;
		15'h047a: char_row_bitmap <= 16'b0011000000110000;
		15'h047b: char_row_bitmap <= 16'b0011100001110000;
		15'h047c: char_row_bitmap <= 16'b0001111111110000;
		15'h047d: char_row_bitmap <= 16'b0000111110110000;
		15'h047e: char_row_bitmap <= 16'b0000000000110000;
		15'h047f: char_row_bitmap <= 16'b0000000000110000;
		15'h0480: char_row_bitmap <= 16'b0000000000110000;
		15'h0481: char_row_bitmap <= 16'b0000000001110000;
		15'h0482: char_row_bitmap <= 16'b0000111111100000;
		15'h0483: char_row_bitmap <= 16'b0000111111000000;
		15'h0484: char_row_bitmap <= 16'b0000000000000000;
		15'h0485: char_row_bitmap <= 16'b0000000000000000;
		15'h0486: char_row_bitmap <= 16'b0000000000000000;
		15'h0487: char_row_bitmap <= 16'b0000000000000000;
		15'h0488: char_row_bitmap <= 16'b0000000000000000;
		15'h0489: char_row_bitmap <= 16'b0000000000000000;
		15'h048a: char_row_bitmap <= 16'b0000000000000000;
		15'h048b: char_row_bitmap <= 16'b0000000000000000;
		15'h048c: char_row_bitmap <= 16'b0000000000000000;
		15'h048d: char_row_bitmap <= 16'b0000000000000000;
		15'h048e: char_row_bitmap <= 16'b0000110000000000;
		15'h048f: char_row_bitmap <= 16'b0000110000000000;
		15'h0490: char_row_bitmap <= 16'b0000000000000000;
		15'h0491: char_row_bitmap <= 16'b0000000000000000;
		15'h0492: char_row_bitmap <= 16'b0000000000000000;
		15'h0493: char_row_bitmap <= 16'b0000000000000000;
		15'h0494: char_row_bitmap <= 16'b0000000000000000;
		15'h0495: char_row_bitmap <= 16'b0000000000000000;
		15'h0496: char_row_bitmap <= 16'b0000110000000000;
		15'h0497: char_row_bitmap <= 16'b0000110000000000;
		15'h0498: char_row_bitmap <= 16'b0000000000000000;
		15'h0499: char_row_bitmap <= 16'b0000000000000000;
		15'h049a: char_row_bitmap <= 16'b0000000000000000;
		15'h049b: char_row_bitmap <= 16'b0000000000000000;
		15'h049c: char_row_bitmap <= 16'b0000000000000000;
		15'h049d: char_row_bitmap <= 16'b0000000000000000;
		15'h049e: char_row_bitmap <= 16'b0000000000000000;
		15'h049f: char_row_bitmap <= 16'b0000000000000000;
		15'h04a0: char_row_bitmap <= 16'b0000000000000000;
		15'h04a1: char_row_bitmap <= 16'b0000000000000000;
		15'h04a2: char_row_bitmap <= 16'b0000110000000000;
		15'h04a3: char_row_bitmap <= 16'b0000110000000000;
		15'h04a4: char_row_bitmap <= 16'b0000000000000000;
		15'h04a5: char_row_bitmap <= 16'b0000000000000000;
		15'h04a6: char_row_bitmap <= 16'b0000000000000000;
		15'h04a7: char_row_bitmap <= 16'b0000000000000000;
		15'h04a8: char_row_bitmap <= 16'b0000110000000000;
		15'h04a9: char_row_bitmap <= 16'b0000110000000000;
		15'h04aa: char_row_bitmap <= 16'b0000110000000000;
		15'h04ab: char_row_bitmap <= 16'b0001110000000000;
		15'h04ac: char_row_bitmap <= 16'b0011100000000000;
		15'h04ad: char_row_bitmap <= 16'b0011000000000000;
		15'h04ae: char_row_bitmap <= 16'b0000000000000000;
		15'h04af: char_row_bitmap <= 16'b0000000000000000;
		15'h04b0: char_row_bitmap <= 16'b0000000000000000;
		15'h04b1: char_row_bitmap <= 16'b0000000000000000;
		15'h04b2: char_row_bitmap <= 16'b0000000000110000;
		15'h04b3: char_row_bitmap <= 16'b0000000001110000;
		15'h04b4: char_row_bitmap <= 16'b0000000011100000;
		15'h04b5: char_row_bitmap <= 16'b0000000111000000;
		15'h04b6: char_row_bitmap <= 16'b0000001110000000;
		15'h04b7: char_row_bitmap <= 16'b0000011100000000;
		15'h04b8: char_row_bitmap <= 16'b0000111000000000;
		15'h04b9: char_row_bitmap <= 16'b0001110000000000;
		15'h04ba: char_row_bitmap <= 16'b0000111000000000;
		15'h04bb: char_row_bitmap <= 16'b0000011100000000;
		15'h04bc: char_row_bitmap <= 16'b0000001110000000;
		15'h04bd: char_row_bitmap <= 16'b0000000111000000;
		15'h04be: char_row_bitmap <= 16'b0000000011100000;
		15'h04bf: char_row_bitmap <= 16'b0000000001110000;
		15'h04c0: char_row_bitmap <= 16'b0000000000110000;
		15'h04c1: char_row_bitmap <= 16'b0000000000000000;
		15'h04c2: char_row_bitmap <= 16'b0000000000000000;
		15'h04c3: char_row_bitmap <= 16'b0000000000000000;
		15'h04c4: char_row_bitmap <= 16'b0000000000000000;
		15'h04c5: char_row_bitmap <= 16'b0000000000000000;
		15'h04c6: char_row_bitmap <= 16'b0000000000000000;
		15'h04c7: char_row_bitmap <= 16'b0000000000000000;
		15'h04c8: char_row_bitmap <= 16'b0000000000000000;
		15'h04c9: char_row_bitmap <= 16'b0000000000000000;
		15'h04ca: char_row_bitmap <= 16'b0011111111110000;
		15'h04cb: char_row_bitmap <= 16'b0011111111110000;
		15'h04cc: char_row_bitmap <= 16'b0000000000000000;
		15'h04cd: char_row_bitmap <= 16'b0000000000000000;
		15'h04ce: char_row_bitmap <= 16'b0011111111110000;
		15'h04cf: char_row_bitmap <= 16'b0011111111110000;
		15'h04d0: char_row_bitmap <= 16'b0000000000000000;
		15'h04d1: char_row_bitmap <= 16'b0000000000000000;
		15'h04d2: char_row_bitmap <= 16'b0000000000000000;
		15'h04d3: char_row_bitmap <= 16'b0000000000000000;
		15'h04d4: char_row_bitmap <= 16'b0000000000000000;
		15'h04d5: char_row_bitmap <= 16'b0000000000000000;
		15'h04d6: char_row_bitmap <= 16'b0000000000000000;
		15'h04d7: char_row_bitmap <= 16'b0000000000000000;
		15'h04d8: char_row_bitmap <= 16'b0000000000000000;
		15'h04d9: char_row_bitmap <= 16'b0000000000000000;
		15'h04da: char_row_bitmap <= 16'b0011000000000000;
		15'h04db: char_row_bitmap <= 16'b0011100000000000;
		15'h04dc: char_row_bitmap <= 16'b0001110000000000;
		15'h04dd: char_row_bitmap <= 16'b0000111000000000;
		15'h04de: char_row_bitmap <= 16'b0000011100000000;
		15'h04df: char_row_bitmap <= 16'b0000001110000000;
		15'h04e0: char_row_bitmap <= 16'b0000000111000000;
		15'h04e1: char_row_bitmap <= 16'b0000000011100000;
		15'h04e2: char_row_bitmap <= 16'b0000000111000000;
		15'h04e3: char_row_bitmap <= 16'b0000001110000000;
		15'h04e4: char_row_bitmap <= 16'b0000011100000000;
		15'h04e5: char_row_bitmap <= 16'b0000111000000000;
		15'h04e6: char_row_bitmap <= 16'b0001110000000000;
		15'h04e7: char_row_bitmap <= 16'b0011100000000000;
		15'h04e8: char_row_bitmap <= 16'b0011000000000000;
		15'h04e9: char_row_bitmap <= 16'b0000000000000000;
		15'h04ea: char_row_bitmap <= 16'b0000000000000000;
		15'h04eb: char_row_bitmap <= 16'b0000000000000000;
		15'h04ec: char_row_bitmap <= 16'b0000000000000000;
		15'h04ed: char_row_bitmap <= 16'b0000000000000000;
		15'h04ee: char_row_bitmap <= 16'b0000111111000000;
		15'h04ef: char_row_bitmap <= 16'b0001111111100000;
		15'h04f0: char_row_bitmap <= 16'b0011100001110000;
		15'h04f1: char_row_bitmap <= 16'b0011000000110000;
		15'h04f2: char_row_bitmap <= 16'b0000000000110000;
		15'h04f3: char_row_bitmap <= 16'b0000000001110000;
		15'h04f4: char_row_bitmap <= 16'b0000000011100000;
		15'h04f5: char_row_bitmap <= 16'b0000000111000000;
		15'h04f6: char_row_bitmap <= 16'b0000001110000000;
		15'h04f7: char_row_bitmap <= 16'b0000001100000000;
		15'h04f8: char_row_bitmap <= 16'b0000000000000000;
		15'h04f9: char_row_bitmap <= 16'b0000000000000000;
		15'h04fa: char_row_bitmap <= 16'b0000001100000000;
		15'h04fb: char_row_bitmap <= 16'b0000001100000000;
		15'h04fc: char_row_bitmap <= 16'b0000000000000000;
		15'h04fd: char_row_bitmap <= 16'b0000000000000000;
		15'h04fe: char_row_bitmap <= 16'b0000000000000000;
		15'h04ff: char_row_bitmap <= 16'b0000000000000000;
		15'h0500: char_row_bitmap <= 16'b0000000000000000;
		15'h0501: char_row_bitmap <= 16'b0000000000000000;
		15'h0502: char_row_bitmap <= 16'b0000111111000000;
		15'h0503: char_row_bitmap <= 16'b0001111111100000;
		15'h0504: char_row_bitmap <= 16'b0011100001110000;
		15'h0505: char_row_bitmap <= 16'b0011000000110000;
		15'h0506: char_row_bitmap <= 16'b0011000111110000;
		15'h0507: char_row_bitmap <= 16'b0011001111110000;
		15'h0508: char_row_bitmap <= 16'b0011001100110000;
		15'h0509: char_row_bitmap <= 16'b0011001100110000;
		15'h050a: char_row_bitmap <= 16'b0011001111110000;
		15'h050b: char_row_bitmap <= 16'b0011000111100000;
		15'h050c: char_row_bitmap <= 16'b0011000000000000;
		15'h050d: char_row_bitmap <= 16'b0011100000000000;
		15'h050e: char_row_bitmap <= 16'b0001111111000000;
		15'h050f: char_row_bitmap <= 16'b0000111111000000;
		15'h0510: char_row_bitmap <= 16'b0000000000000000;
		15'h0511: char_row_bitmap <= 16'b0000000000000000;
		15'h0512: char_row_bitmap <= 16'b0000000000000000;
		15'h0513: char_row_bitmap <= 16'b0000000000000000;
		15'h0514: char_row_bitmap <= 16'b0000000000000000;
		15'h0515: char_row_bitmap <= 16'b0000000000000000;
		15'h0516: char_row_bitmap <= 16'b0000111111000000;
		15'h0517: char_row_bitmap <= 16'b0001111111100000;
		15'h0518: char_row_bitmap <= 16'b0011100001110000;
		15'h0519: char_row_bitmap <= 16'b0011000000110000;
		15'h051a: char_row_bitmap <= 16'b0011000000110000;
		15'h051b: char_row_bitmap <= 16'b0011000000110000;
		15'h051c: char_row_bitmap <= 16'b0011000000110000;
		15'h051d: char_row_bitmap <= 16'b0011000000110000;
		15'h051e: char_row_bitmap <= 16'b0011111111110000;
		15'h051f: char_row_bitmap <= 16'b0011111111110000;
		15'h0520: char_row_bitmap <= 16'b0011000000110000;
		15'h0521: char_row_bitmap <= 16'b0011000000110000;
		15'h0522: char_row_bitmap <= 16'b0011000000110000;
		15'h0523: char_row_bitmap <= 16'b0011000000110000;
		15'h0524: char_row_bitmap <= 16'b0000000000000000;
		15'h0525: char_row_bitmap <= 16'b0000000000000000;
		15'h0526: char_row_bitmap <= 16'b0000000000000000;
		15'h0527: char_row_bitmap <= 16'b0000000000000000;
		15'h0528: char_row_bitmap <= 16'b0000000000000000;
		15'h0529: char_row_bitmap <= 16'b0000000000000000;
		15'h052a: char_row_bitmap <= 16'b0011111111000000;
		15'h052b: char_row_bitmap <= 16'b0011111111100000;
		15'h052c: char_row_bitmap <= 16'b0011000001110000;
		15'h052d: char_row_bitmap <= 16'b0011000000110000;
		15'h052e: char_row_bitmap <= 16'b0011000000110000;
		15'h052f: char_row_bitmap <= 16'b0011000001110000;
		15'h0530: char_row_bitmap <= 16'b0011111111100000;
		15'h0531: char_row_bitmap <= 16'b0011111111100000;
		15'h0532: char_row_bitmap <= 16'b0011000001110000;
		15'h0533: char_row_bitmap <= 16'b0011000000110000;
		15'h0534: char_row_bitmap <= 16'b0011000000110000;
		15'h0535: char_row_bitmap <= 16'b0011000001110000;
		15'h0536: char_row_bitmap <= 16'b0011111111100000;
		15'h0537: char_row_bitmap <= 16'b0011111111000000;
		15'h0538: char_row_bitmap <= 16'b0000000000000000;
		15'h0539: char_row_bitmap <= 16'b0000000000000000;
		15'h053a: char_row_bitmap <= 16'b0000000000000000;
		15'h053b: char_row_bitmap <= 16'b0000000000000000;
		15'h053c: char_row_bitmap <= 16'b0000000000000000;
		15'h053d: char_row_bitmap <= 16'b0000000000000000;
		15'h053e: char_row_bitmap <= 16'b0000111111000000;
		15'h053f: char_row_bitmap <= 16'b0001111111100000;
		15'h0540: char_row_bitmap <= 16'b0011100001110000;
		15'h0541: char_row_bitmap <= 16'b0011000000110000;
		15'h0542: char_row_bitmap <= 16'b0011000000000000;
		15'h0543: char_row_bitmap <= 16'b0011000000000000;
		15'h0544: char_row_bitmap <= 16'b0011000000000000;
		15'h0545: char_row_bitmap <= 16'b0011000000000000;
		15'h0546: char_row_bitmap <= 16'b0011000000000000;
		15'h0547: char_row_bitmap <= 16'b0011000000000000;
		15'h0548: char_row_bitmap <= 16'b0011000000110000;
		15'h0549: char_row_bitmap <= 16'b0011100001110000;
		15'h054a: char_row_bitmap <= 16'b0001111111100000;
		15'h054b: char_row_bitmap <= 16'b0000111111000000;
		15'h054c: char_row_bitmap <= 16'b0000000000000000;
		15'h054d: char_row_bitmap <= 16'b0000000000000000;
		15'h054e: char_row_bitmap <= 16'b0000000000000000;
		15'h054f: char_row_bitmap <= 16'b0000000000000000;
		15'h0550: char_row_bitmap <= 16'b0000000000000000;
		15'h0551: char_row_bitmap <= 16'b0000000000000000;
		15'h0552: char_row_bitmap <= 16'b0011111111000000;
		15'h0553: char_row_bitmap <= 16'b0011111111100000;
		15'h0554: char_row_bitmap <= 16'b0011000001110000;
		15'h0555: char_row_bitmap <= 16'b0011000000110000;
		15'h0556: char_row_bitmap <= 16'b0011000000110000;
		15'h0557: char_row_bitmap <= 16'b0011000000110000;
		15'h0558: char_row_bitmap <= 16'b0011000000110000;
		15'h0559: char_row_bitmap <= 16'b0011000000110000;
		15'h055a: char_row_bitmap <= 16'b0011000000110000;
		15'h055b: char_row_bitmap <= 16'b0011000000110000;
		15'h055c: char_row_bitmap <= 16'b0011000000110000;
		15'h055d: char_row_bitmap <= 16'b0011000001110000;
		15'h055e: char_row_bitmap <= 16'b0011111111100000;
		15'h055f: char_row_bitmap <= 16'b0011111111000000;
		15'h0560: char_row_bitmap <= 16'b0000000000000000;
		15'h0561: char_row_bitmap <= 16'b0000000000000000;
		15'h0562: char_row_bitmap <= 16'b0000000000000000;
		15'h0563: char_row_bitmap <= 16'b0000000000000000;
		15'h0564: char_row_bitmap <= 16'b0000000000000000;
		15'h0565: char_row_bitmap <= 16'b0000000000000000;
		15'h0566: char_row_bitmap <= 16'b0011111111110000;
		15'h0567: char_row_bitmap <= 16'b0011111111110000;
		15'h0568: char_row_bitmap <= 16'b0011000000000000;
		15'h0569: char_row_bitmap <= 16'b0011000000000000;
		15'h056a: char_row_bitmap <= 16'b0011000000000000;
		15'h056b: char_row_bitmap <= 16'b0011000000000000;
		15'h056c: char_row_bitmap <= 16'b0011111100000000;
		15'h056d: char_row_bitmap <= 16'b0011111100000000;
		15'h056e: char_row_bitmap <= 16'b0011000000000000;
		15'h056f: char_row_bitmap <= 16'b0011000000000000;
		15'h0570: char_row_bitmap <= 16'b0011000000000000;
		15'h0571: char_row_bitmap <= 16'b0011000000000000;
		15'h0572: char_row_bitmap <= 16'b0011111111110000;
		15'h0573: char_row_bitmap <= 16'b0011111111110000;
		15'h0574: char_row_bitmap <= 16'b0000000000000000;
		15'h0575: char_row_bitmap <= 16'b0000000000000000;
		15'h0576: char_row_bitmap <= 16'b0000000000000000;
		15'h0577: char_row_bitmap <= 16'b0000000000000000;
		15'h0578: char_row_bitmap <= 16'b0000000000000000;
		15'h0579: char_row_bitmap <= 16'b0000000000000000;
		15'h057a: char_row_bitmap <= 16'b0011111111110000;
		15'h057b: char_row_bitmap <= 16'b0011111111110000;
		15'h057c: char_row_bitmap <= 16'b0011000000000000;
		15'h057d: char_row_bitmap <= 16'b0011000000000000;
		15'h057e: char_row_bitmap <= 16'b0011000000000000;
		15'h057f: char_row_bitmap <= 16'b0011000000000000;
		15'h0580: char_row_bitmap <= 16'b0011111100000000;
		15'h0581: char_row_bitmap <= 16'b0011111100000000;
		15'h0582: char_row_bitmap <= 16'b0011000000000000;
		15'h0583: char_row_bitmap <= 16'b0011000000000000;
		15'h0584: char_row_bitmap <= 16'b0011000000000000;
		15'h0585: char_row_bitmap <= 16'b0011000000000000;
		15'h0586: char_row_bitmap <= 16'b0011000000000000;
		15'h0587: char_row_bitmap <= 16'b0011000000000000;
		15'h0588: char_row_bitmap <= 16'b0000000000000000;
		15'h0589: char_row_bitmap <= 16'b0000000000000000;
		15'h058a: char_row_bitmap <= 16'b0000000000000000;
		15'h058b: char_row_bitmap <= 16'b0000000000000000;
		15'h058c: char_row_bitmap <= 16'b0000000000000000;
		15'h058d: char_row_bitmap <= 16'b0000000000000000;
		15'h058e: char_row_bitmap <= 16'b0000111111000000;
		15'h058f: char_row_bitmap <= 16'b0001111111100000;
		15'h0590: char_row_bitmap <= 16'b0011100001110000;
		15'h0591: char_row_bitmap <= 16'b0011000000110000;
		15'h0592: char_row_bitmap <= 16'b0011000000000000;
		15'h0593: char_row_bitmap <= 16'b0011000000000000;
		15'h0594: char_row_bitmap <= 16'b0011000000000000;
		15'h0595: char_row_bitmap <= 16'b0011000000000000;
		15'h0596: char_row_bitmap <= 16'b0011000011110000;
		15'h0597: char_row_bitmap <= 16'b0011000011110000;
		15'h0598: char_row_bitmap <= 16'b0011000000110000;
		15'h0599: char_row_bitmap <= 16'b0011100000110000;
		15'h059a: char_row_bitmap <= 16'b0001111111110000;
		15'h059b: char_row_bitmap <= 16'b0000111111100000;
		15'h059c: char_row_bitmap <= 16'b0000000000000000;
		15'h059d: char_row_bitmap <= 16'b0000000000000000;
		15'h059e: char_row_bitmap <= 16'b0000000000000000;
		15'h059f: char_row_bitmap <= 16'b0000000000000000;
		15'h05a0: char_row_bitmap <= 16'b0000000000000000;
		15'h05a1: char_row_bitmap <= 16'b0000000000000000;
		15'h05a2: char_row_bitmap <= 16'b0011000000110000;
		15'h05a3: char_row_bitmap <= 16'b0011000000110000;
		15'h05a4: char_row_bitmap <= 16'b0011000000110000;
		15'h05a5: char_row_bitmap <= 16'b0011000000110000;
		15'h05a6: char_row_bitmap <= 16'b0011000000110000;
		15'h05a7: char_row_bitmap <= 16'b0011000000110000;
		15'h05a8: char_row_bitmap <= 16'b0011111111110000;
		15'h05a9: char_row_bitmap <= 16'b0011111111110000;
		15'h05aa: char_row_bitmap <= 16'b0011000000110000;
		15'h05ab: char_row_bitmap <= 16'b0011000000110000;
		15'h05ac: char_row_bitmap <= 16'b0011000000110000;
		15'h05ad: char_row_bitmap <= 16'b0011000000110000;
		15'h05ae: char_row_bitmap <= 16'b0011000000110000;
		15'h05af: char_row_bitmap <= 16'b0011000000110000;
		15'h05b0: char_row_bitmap <= 16'b0000000000000000;
		15'h05b1: char_row_bitmap <= 16'b0000000000000000;
		15'h05b2: char_row_bitmap <= 16'b0000000000000000;
		15'h05b3: char_row_bitmap <= 16'b0000000000000000;
		15'h05b4: char_row_bitmap <= 16'b0000000000000000;
		15'h05b5: char_row_bitmap <= 16'b0000000000000000;
		15'h05b6: char_row_bitmap <= 16'b0000111111000000;
		15'h05b7: char_row_bitmap <= 16'b0000111111000000;
		15'h05b8: char_row_bitmap <= 16'b0000001100000000;
		15'h05b9: char_row_bitmap <= 16'b0000001100000000;
		15'h05ba: char_row_bitmap <= 16'b0000001100000000;
		15'h05bb: char_row_bitmap <= 16'b0000001100000000;
		15'h05bc: char_row_bitmap <= 16'b0000001100000000;
		15'h05bd: char_row_bitmap <= 16'b0000001100000000;
		15'h05be: char_row_bitmap <= 16'b0000001100000000;
		15'h05bf: char_row_bitmap <= 16'b0000001100000000;
		15'h05c0: char_row_bitmap <= 16'b0000001100000000;
		15'h05c1: char_row_bitmap <= 16'b0000001100000000;
		15'h05c2: char_row_bitmap <= 16'b0000111111000000;
		15'h05c3: char_row_bitmap <= 16'b0000111111000000;
		15'h05c4: char_row_bitmap <= 16'b0000000000000000;
		15'h05c5: char_row_bitmap <= 16'b0000000000000000;
		15'h05c6: char_row_bitmap <= 16'b0000000000000000;
		15'h05c7: char_row_bitmap <= 16'b0000000000000000;
		15'h05c8: char_row_bitmap <= 16'b0000000000000000;
		15'h05c9: char_row_bitmap <= 16'b0000000000000000;
		15'h05ca: char_row_bitmap <= 16'b0000001111110000;
		15'h05cb: char_row_bitmap <= 16'b0000001111110000;
		15'h05cc: char_row_bitmap <= 16'b0000000011000000;
		15'h05cd: char_row_bitmap <= 16'b0000000011000000;
		15'h05ce: char_row_bitmap <= 16'b0000000011000000;
		15'h05cf: char_row_bitmap <= 16'b0000000011000000;
		15'h05d0: char_row_bitmap <= 16'b0000000011000000;
		15'h05d1: char_row_bitmap <= 16'b0000000011000000;
		15'h05d2: char_row_bitmap <= 16'b0000000011000000;
		15'h05d3: char_row_bitmap <= 16'b0000000011000000;
		15'h05d4: char_row_bitmap <= 16'b0011000011000000;
		15'h05d5: char_row_bitmap <= 16'b0011100111000000;
		15'h05d6: char_row_bitmap <= 16'b0001111110000000;
		15'h05d7: char_row_bitmap <= 16'b0000111100000000;
		15'h05d8: char_row_bitmap <= 16'b0000000000000000;
		15'h05d9: char_row_bitmap <= 16'b0000000000000000;
		15'h05da: char_row_bitmap <= 16'b0000000000000000;
		15'h05db: char_row_bitmap <= 16'b0000000000000000;
		15'h05dc: char_row_bitmap <= 16'b0000000000000000;
		15'h05dd: char_row_bitmap <= 16'b0000000000000000;
		15'h05de: char_row_bitmap <= 16'b0011000000110000;
		15'h05df: char_row_bitmap <= 16'b0011000001110000;
		15'h05e0: char_row_bitmap <= 16'b0011000011100000;
		15'h05e1: char_row_bitmap <= 16'b0011000111000000;
		15'h05e2: char_row_bitmap <= 16'b0011001110000000;
		15'h05e3: char_row_bitmap <= 16'b0011011100000000;
		15'h05e4: char_row_bitmap <= 16'b0011111000000000;
		15'h05e5: char_row_bitmap <= 16'b0011111000000000;
		15'h05e6: char_row_bitmap <= 16'b0011011100000000;
		15'h05e7: char_row_bitmap <= 16'b0011001110000000;
		15'h05e8: char_row_bitmap <= 16'b0011000111000000;
		15'h05e9: char_row_bitmap <= 16'b0011000011100000;
		15'h05ea: char_row_bitmap <= 16'b0011000001110000;
		15'h05eb: char_row_bitmap <= 16'b0011000000110000;
		15'h05ec: char_row_bitmap <= 16'b0000000000000000;
		15'h05ed: char_row_bitmap <= 16'b0000000000000000;
		15'h05ee: char_row_bitmap <= 16'b0000000000000000;
		15'h05ef: char_row_bitmap <= 16'b0000000000000000;
		15'h05f0: char_row_bitmap <= 16'b0000000000000000;
		15'h05f1: char_row_bitmap <= 16'b0000000000000000;
		15'h05f2: char_row_bitmap <= 16'b0011000000000000;
		15'h05f3: char_row_bitmap <= 16'b0011000000000000;
		15'h05f4: char_row_bitmap <= 16'b0011000000000000;
		15'h05f5: char_row_bitmap <= 16'b0011000000000000;
		15'h05f6: char_row_bitmap <= 16'b0011000000000000;
		15'h05f7: char_row_bitmap <= 16'b0011000000000000;
		15'h05f8: char_row_bitmap <= 16'b0011000000000000;
		15'h05f9: char_row_bitmap <= 16'b0011000000000000;
		15'h05fa: char_row_bitmap <= 16'b0011000000000000;
		15'h05fb: char_row_bitmap <= 16'b0011000000000000;
		15'h05fc: char_row_bitmap <= 16'b0011000000000000;
		15'h05fd: char_row_bitmap <= 16'b0011000000000000;
		15'h05fe: char_row_bitmap <= 16'b0011111111110000;
		15'h05ff: char_row_bitmap <= 16'b0011111111110000;
		15'h0600: char_row_bitmap <= 16'b0000000000000000;
		15'h0601: char_row_bitmap <= 16'b0000000000000000;
		15'h0602: char_row_bitmap <= 16'b0000000000000000;
		15'h0603: char_row_bitmap <= 16'b0000000000000000;
		15'h0604: char_row_bitmap <= 16'b0000000000000000;
		15'h0605: char_row_bitmap <= 16'b0000000000000000;
		15'h0606: char_row_bitmap <= 16'b0011000000110000;
		15'h0607: char_row_bitmap <= 16'b0011100001110000;
		15'h0608: char_row_bitmap <= 16'b0011110011110000;
		15'h0609: char_row_bitmap <= 16'b0011111111110000;
		15'h060a: char_row_bitmap <= 16'b0011011110110000;
		15'h060b: char_row_bitmap <= 16'b0011001100110000;
		15'h060c: char_row_bitmap <= 16'b0011001100110000;
		15'h060d: char_row_bitmap <= 16'b0011000000110000;
		15'h060e: char_row_bitmap <= 16'b0011000000110000;
		15'h060f: char_row_bitmap <= 16'b0011000000110000;
		15'h0610: char_row_bitmap <= 16'b0011000000110000;
		15'h0611: char_row_bitmap <= 16'b0011000000110000;
		15'h0612: char_row_bitmap <= 16'b0011000000110000;
		15'h0613: char_row_bitmap <= 16'b0011000000110000;
		15'h0614: char_row_bitmap <= 16'b0000000000000000;
		15'h0615: char_row_bitmap <= 16'b0000000000000000;
		15'h0616: char_row_bitmap <= 16'b0000000000000000;
		15'h0617: char_row_bitmap <= 16'b0000000000000000;
		15'h0618: char_row_bitmap <= 16'b0000000000000000;
		15'h0619: char_row_bitmap <= 16'b0000000000000000;
		15'h061a: char_row_bitmap <= 16'b0011000000110000;
		15'h061b: char_row_bitmap <= 16'b0011000000110000;
		15'h061c: char_row_bitmap <= 16'b0011000000110000;
		15'h061d: char_row_bitmap <= 16'b0011100000110000;
		15'h061e: char_row_bitmap <= 16'b0011110000110000;
		15'h061f: char_row_bitmap <= 16'b0011111000110000;
		15'h0620: char_row_bitmap <= 16'b0011011100110000;
		15'h0621: char_row_bitmap <= 16'b0011001110110000;
		15'h0622: char_row_bitmap <= 16'b0011000111110000;
		15'h0623: char_row_bitmap <= 16'b0011000011110000;
		15'h0624: char_row_bitmap <= 16'b0011000001110000;
		15'h0625: char_row_bitmap <= 16'b0011000000110000;
		15'h0626: char_row_bitmap <= 16'b0011000000110000;
		15'h0627: char_row_bitmap <= 16'b0011000000110000;
		15'h0628: char_row_bitmap <= 16'b0000000000000000;
		15'h0629: char_row_bitmap <= 16'b0000000000000000;
		15'h062a: char_row_bitmap <= 16'b0000000000000000;
		15'h062b: char_row_bitmap <= 16'b0000000000000000;
		15'h062c: char_row_bitmap <= 16'b0000000000000000;
		15'h062d: char_row_bitmap <= 16'b0000000000000000;
		15'h062e: char_row_bitmap <= 16'b0000111111000000;
		15'h062f: char_row_bitmap <= 16'b0001111111100000;
		15'h0630: char_row_bitmap <= 16'b0011100001110000;
		15'h0631: char_row_bitmap <= 16'b0011000000110000;
		15'h0632: char_row_bitmap <= 16'b0011000000110000;
		15'h0633: char_row_bitmap <= 16'b0011000000110000;
		15'h0634: char_row_bitmap <= 16'b0011000000110000;
		15'h0635: char_row_bitmap <= 16'b0011000000110000;
		15'h0636: char_row_bitmap <= 16'b0011000000110000;
		15'h0637: char_row_bitmap <= 16'b0011000000110000;
		15'h0638: char_row_bitmap <= 16'b0011000000110000;
		15'h0639: char_row_bitmap <= 16'b0011100001110000;
		15'h063a: char_row_bitmap <= 16'b0001111111100000;
		15'h063b: char_row_bitmap <= 16'b0000111111000000;
		15'h063c: char_row_bitmap <= 16'b0000000000000000;
		15'h063d: char_row_bitmap <= 16'b0000000000000000;
		15'h063e: char_row_bitmap <= 16'b0000000000000000;
		15'h063f: char_row_bitmap <= 16'b0000000000000000;
		15'h0640: char_row_bitmap <= 16'b0000000000000000;
		15'h0641: char_row_bitmap <= 16'b0000000000000000;
		15'h0642: char_row_bitmap <= 16'b0011111111000000;
		15'h0643: char_row_bitmap <= 16'b0011111111100000;
		15'h0644: char_row_bitmap <= 16'b0011000001110000;
		15'h0645: char_row_bitmap <= 16'b0011000000110000;
		15'h0646: char_row_bitmap <= 16'b0011000000110000;
		15'h0647: char_row_bitmap <= 16'b0011000001110000;
		15'h0648: char_row_bitmap <= 16'b0011111111100000;
		15'h0649: char_row_bitmap <= 16'b0011111111000000;
		15'h064a: char_row_bitmap <= 16'b0011000000000000;
		15'h064b: char_row_bitmap <= 16'b0011000000000000;
		15'h064c: char_row_bitmap <= 16'b0011000000000000;
		15'h064d: char_row_bitmap <= 16'b0011000000000000;
		15'h064e: char_row_bitmap <= 16'b0011000000000000;
		15'h064f: char_row_bitmap <= 16'b0011000000000000;
		15'h0650: char_row_bitmap <= 16'b0000000000000000;
		15'h0651: char_row_bitmap <= 16'b0000000000000000;
		15'h0652: char_row_bitmap <= 16'b0000000000000000;
		15'h0653: char_row_bitmap <= 16'b0000000000000000;
		15'h0654: char_row_bitmap <= 16'b0000000000000000;
		15'h0655: char_row_bitmap <= 16'b0000000000000000;
		15'h0656: char_row_bitmap <= 16'b0000111111000000;
		15'h0657: char_row_bitmap <= 16'b0001111111100000;
		15'h0658: char_row_bitmap <= 16'b0011100001110000;
		15'h0659: char_row_bitmap <= 16'b0011000000110000;
		15'h065a: char_row_bitmap <= 16'b0011000000110000;
		15'h065b: char_row_bitmap <= 16'b0011000000110000;
		15'h065c: char_row_bitmap <= 16'b0011000000110000;
		15'h065d: char_row_bitmap <= 16'b0011000000110000;
		15'h065e: char_row_bitmap <= 16'b0011001100110000;
		15'h065f: char_row_bitmap <= 16'b0011001110110000;
		15'h0660: char_row_bitmap <= 16'b0011000111000000;
		15'h0661: char_row_bitmap <= 16'b0011000011100000;
		15'h0662: char_row_bitmap <= 16'b0001111101110000;
		15'h0663: char_row_bitmap <= 16'b0000111100110000;
		15'h0664: char_row_bitmap <= 16'b0000000000000000;
		15'h0665: char_row_bitmap <= 16'b0000000000000000;
		15'h0666: char_row_bitmap <= 16'b0000000000000000;
		15'h0667: char_row_bitmap <= 16'b0000000000000000;
		15'h0668: char_row_bitmap <= 16'b0000000000000000;
		15'h0669: char_row_bitmap <= 16'b0000000000000000;
		15'h066a: char_row_bitmap <= 16'b0011111111000000;
		15'h066b: char_row_bitmap <= 16'b0011111111100000;
		15'h066c: char_row_bitmap <= 16'b0011000001110000;
		15'h066d: char_row_bitmap <= 16'b0011000000110000;
		15'h066e: char_row_bitmap <= 16'b0011000000110000;
		15'h066f: char_row_bitmap <= 16'b0011000001110000;
		15'h0670: char_row_bitmap <= 16'b0011111111100000;
		15'h0671: char_row_bitmap <= 16'b0011111111000000;
		15'h0672: char_row_bitmap <= 16'b0011011100000000;
		15'h0673: char_row_bitmap <= 16'b0011001110000000;
		15'h0674: char_row_bitmap <= 16'b0011000111000000;
		15'h0675: char_row_bitmap <= 16'b0011000011100000;
		15'h0676: char_row_bitmap <= 16'b0011000001110000;
		15'h0677: char_row_bitmap <= 16'b0011000000110000;
		15'h0678: char_row_bitmap <= 16'b0000000000000000;
		15'h0679: char_row_bitmap <= 16'b0000000000000000;
		15'h067a: char_row_bitmap <= 16'b0000000000000000;
		15'h067b: char_row_bitmap <= 16'b0000000000000000;
		15'h067c: char_row_bitmap <= 16'b0000000000000000;
		15'h067d: char_row_bitmap <= 16'b0000000000000000;
		15'h067e: char_row_bitmap <= 16'b0000111111000000;
		15'h067f: char_row_bitmap <= 16'b0001111111100000;
		15'h0680: char_row_bitmap <= 16'b0011100001110000;
		15'h0681: char_row_bitmap <= 16'b0011000000110000;
		15'h0682: char_row_bitmap <= 16'b0011000000000000;
		15'h0683: char_row_bitmap <= 16'b0011100000000000;
		15'h0684: char_row_bitmap <= 16'b0001111111000000;
		15'h0685: char_row_bitmap <= 16'b0000111111100000;
		15'h0686: char_row_bitmap <= 16'b0000000001110000;
		15'h0687: char_row_bitmap <= 16'b0000000000110000;
		15'h0688: char_row_bitmap <= 16'b0011000000110000;
		15'h0689: char_row_bitmap <= 16'b0011100001110000;
		15'h068a: char_row_bitmap <= 16'b0001111111100000;
		15'h068b: char_row_bitmap <= 16'b0000111111000000;
		15'h068c: char_row_bitmap <= 16'b0000000000000000;
		15'h068d: char_row_bitmap <= 16'b0000000000000000;
		15'h068e: char_row_bitmap <= 16'b0000000000000000;
		15'h068f: char_row_bitmap <= 16'b0000000000000000;
		15'h0690: char_row_bitmap <= 16'b0000000000000000;
		15'h0691: char_row_bitmap <= 16'b0000000000000000;
		15'h0692: char_row_bitmap <= 16'b0011111111110000;
		15'h0693: char_row_bitmap <= 16'b0011111111110000;
		15'h0694: char_row_bitmap <= 16'b0000001100000000;
		15'h0695: char_row_bitmap <= 16'b0000001100000000;
		15'h0696: char_row_bitmap <= 16'b0000001100000000;
		15'h0697: char_row_bitmap <= 16'b0000001100000000;
		15'h0698: char_row_bitmap <= 16'b0000001100000000;
		15'h0699: char_row_bitmap <= 16'b0000001100000000;
		15'h069a: char_row_bitmap <= 16'b0000001100000000;
		15'h069b: char_row_bitmap <= 16'b0000001100000000;
		15'h069c: char_row_bitmap <= 16'b0000001100000000;
		15'h069d: char_row_bitmap <= 16'b0000001100000000;
		15'h069e: char_row_bitmap <= 16'b0000001100000000;
		15'h069f: char_row_bitmap <= 16'b0000001100000000;
		15'h06a0: char_row_bitmap <= 16'b0000000000000000;
		15'h06a1: char_row_bitmap <= 16'b0000000000000000;
		15'h06a2: char_row_bitmap <= 16'b0000000000000000;
		15'h06a3: char_row_bitmap <= 16'b0000000000000000;
		15'h06a4: char_row_bitmap <= 16'b0000000000000000;
		15'h06a5: char_row_bitmap <= 16'b0000000000000000;
		15'h06a6: char_row_bitmap <= 16'b0011000000110000;
		15'h06a7: char_row_bitmap <= 16'b0011000000110000;
		15'h06a8: char_row_bitmap <= 16'b0011000000110000;
		15'h06a9: char_row_bitmap <= 16'b0011000000110000;
		15'h06aa: char_row_bitmap <= 16'b0011000000110000;
		15'h06ab: char_row_bitmap <= 16'b0011000000110000;
		15'h06ac: char_row_bitmap <= 16'b0011000000110000;
		15'h06ad: char_row_bitmap <= 16'b0011000000110000;
		15'h06ae: char_row_bitmap <= 16'b0011000000110000;
		15'h06af: char_row_bitmap <= 16'b0011000000110000;
		15'h06b0: char_row_bitmap <= 16'b0011000000110000;
		15'h06b1: char_row_bitmap <= 16'b0011100001110000;
		15'h06b2: char_row_bitmap <= 16'b0001111111100000;
		15'h06b3: char_row_bitmap <= 16'b0000111111000000;
		15'h06b4: char_row_bitmap <= 16'b0000000000000000;
		15'h06b5: char_row_bitmap <= 16'b0000000000000000;
		15'h06b6: char_row_bitmap <= 16'b0000000000000000;
		15'h06b7: char_row_bitmap <= 16'b0000000000000000;
		15'h06b8: char_row_bitmap <= 16'b0000000000000000;
		15'h06b9: char_row_bitmap <= 16'b0000000000000000;
		15'h06ba: char_row_bitmap <= 16'b0011000000110000;
		15'h06bb: char_row_bitmap <= 16'b0011000000110000;
		15'h06bc: char_row_bitmap <= 16'b0011000000110000;
		15'h06bd: char_row_bitmap <= 16'b0011000000110000;
		15'h06be: char_row_bitmap <= 16'b0011000000110000;
		15'h06bf: char_row_bitmap <= 16'b0011100001110000;
		15'h06c0: char_row_bitmap <= 16'b0001100001100000;
		15'h06c1: char_row_bitmap <= 16'b0000110011000000;
		15'h06c2: char_row_bitmap <= 16'b0000110011000000;
		15'h06c3: char_row_bitmap <= 16'b0000110011000000;
		15'h06c4: char_row_bitmap <= 16'b0000011110000000;
		15'h06c5: char_row_bitmap <= 16'b0000011110000000;
		15'h06c6: char_row_bitmap <= 16'b0000001100000000;
		15'h06c7: char_row_bitmap <= 16'b0000001100000000;
		15'h06c8: char_row_bitmap <= 16'b0000000000000000;
		15'h06c9: char_row_bitmap <= 16'b0000000000000000;
		15'h06ca: char_row_bitmap <= 16'b0000000000000000;
		15'h06cb: char_row_bitmap <= 16'b0000000000000000;
		15'h06cc: char_row_bitmap <= 16'b0000000000000000;
		15'h06cd: char_row_bitmap <= 16'b0000000000000000;
		15'h06ce: char_row_bitmap <= 16'b0011000000110000;
		15'h06cf: char_row_bitmap <= 16'b0011000000110000;
		15'h06d0: char_row_bitmap <= 16'b0011000000110000;
		15'h06d1: char_row_bitmap <= 16'b0011000000110000;
		15'h06d2: char_row_bitmap <= 16'b0011000000110000;
		15'h06d3: char_row_bitmap <= 16'b0011000000110000;
		15'h06d4: char_row_bitmap <= 16'b0011001100110000;
		15'h06d5: char_row_bitmap <= 16'b0011001100110000;
		15'h06d6: char_row_bitmap <= 16'b0011001100110000;
		15'h06d7: char_row_bitmap <= 16'b0011001100110000;
		15'h06d8: char_row_bitmap <= 16'b0011001100110000;
		15'h06d9: char_row_bitmap <= 16'b0011111111110000;
		15'h06da: char_row_bitmap <= 16'b0001111111100000;
		15'h06db: char_row_bitmap <= 16'b0000110011000000;
		15'h06dc: char_row_bitmap <= 16'b0000000000000000;
		15'h06dd: char_row_bitmap <= 16'b0000000000000000;
		15'h06de: char_row_bitmap <= 16'b0000000000000000;
		15'h06df: char_row_bitmap <= 16'b0000000000000000;
		15'h06e0: char_row_bitmap <= 16'b0000000000000000;
		15'h06e1: char_row_bitmap <= 16'b0000000000000000;
		15'h06e2: char_row_bitmap <= 16'b0011000000110000;
		15'h06e3: char_row_bitmap <= 16'b0011000000110000;
		15'h06e4: char_row_bitmap <= 16'b0011100001110000;
		15'h06e5: char_row_bitmap <= 16'b0001100001100000;
		15'h06e6: char_row_bitmap <= 16'b0001110011100000;
		15'h06e7: char_row_bitmap <= 16'b0000111111000000;
		15'h06e8: char_row_bitmap <= 16'b0000011110000000;
		15'h06e9: char_row_bitmap <= 16'b0000011110000000;
		15'h06ea: char_row_bitmap <= 16'b0000111111000000;
		15'h06eb: char_row_bitmap <= 16'b0001110011100000;
		15'h06ec: char_row_bitmap <= 16'b0001100001100000;
		15'h06ed: char_row_bitmap <= 16'b0011100001110000;
		15'h06ee: char_row_bitmap <= 16'b0011000000110000;
		15'h06ef: char_row_bitmap <= 16'b0011000000110000;
		15'h06f0: char_row_bitmap <= 16'b0000000000000000;
		15'h06f1: char_row_bitmap <= 16'b0000000000000000;
		15'h06f2: char_row_bitmap <= 16'b0000000000000000;
		15'h06f3: char_row_bitmap <= 16'b0000000000000000;
		15'h06f4: char_row_bitmap <= 16'b0000000000000000;
		15'h06f5: char_row_bitmap <= 16'b0000000000000000;
		15'h06f6: char_row_bitmap <= 16'b0011000000110000;
		15'h06f7: char_row_bitmap <= 16'b0011000000110000;
		15'h06f8: char_row_bitmap <= 16'b0011100001110000;
		15'h06f9: char_row_bitmap <= 16'b0001100001100000;
		15'h06fa: char_row_bitmap <= 16'b0001110011100000;
		15'h06fb: char_row_bitmap <= 16'b0000110011000000;
		15'h06fc: char_row_bitmap <= 16'b0000011110000000;
		15'h06fd: char_row_bitmap <= 16'b0000011110000000;
		15'h06fe: char_row_bitmap <= 16'b0000001100000000;
		15'h06ff: char_row_bitmap <= 16'b0000001100000000;
		15'h0700: char_row_bitmap <= 16'b0000001100000000;
		15'h0701: char_row_bitmap <= 16'b0000001100000000;
		15'h0702: char_row_bitmap <= 16'b0000001100000000;
		15'h0703: char_row_bitmap <= 16'b0000001100000000;
		15'h0704: char_row_bitmap <= 16'b0000000000000000;
		15'h0705: char_row_bitmap <= 16'b0000000000000000;
		15'h0706: char_row_bitmap <= 16'b0000000000000000;
		15'h0707: char_row_bitmap <= 16'b0000000000000000;
		15'h0708: char_row_bitmap <= 16'b0000000000000000;
		15'h0709: char_row_bitmap <= 16'b0000000000000000;
		15'h070a: char_row_bitmap <= 16'b0011111111110000;
		15'h070b: char_row_bitmap <= 16'b0011111111110000;
		15'h070c: char_row_bitmap <= 16'b0000000000110000;
		15'h070d: char_row_bitmap <= 16'b0000000001110000;
		15'h070e: char_row_bitmap <= 16'b0000000011100000;
		15'h070f: char_row_bitmap <= 16'b0000000111000000;
		15'h0710: char_row_bitmap <= 16'b0000001110000000;
		15'h0711: char_row_bitmap <= 16'b0000011100000000;
		15'h0712: char_row_bitmap <= 16'b0000111000000000;
		15'h0713: char_row_bitmap <= 16'b0001110000000000;
		15'h0714: char_row_bitmap <= 16'b0011100000000000;
		15'h0715: char_row_bitmap <= 16'b0011000000000000;
		15'h0716: char_row_bitmap <= 16'b0011111111110000;
		15'h0717: char_row_bitmap <= 16'b0011111111110000;
		15'h0718: char_row_bitmap <= 16'b0000000000000000;
		15'h0719: char_row_bitmap <= 16'b0000000000000000;
		15'h071a: char_row_bitmap <= 16'b0000000000000000;
		15'h071b: char_row_bitmap <= 16'b0000000000000000;
		15'h071c: char_row_bitmap <= 16'b0000000000000000;
		15'h071d: char_row_bitmap <= 16'b0000000000000000;
		15'h071e: char_row_bitmap <= 16'b0000001111110000;
		15'h071f: char_row_bitmap <= 16'b0000001111110000;
		15'h0720: char_row_bitmap <= 16'b0000001100000000;
		15'h0721: char_row_bitmap <= 16'b0000001100000000;
		15'h0722: char_row_bitmap <= 16'b0000001100000000;
		15'h0723: char_row_bitmap <= 16'b0000001100000000;
		15'h0724: char_row_bitmap <= 16'b0000001100000000;
		15'h0725: char_row_bitmap <= 16'b0000001100000000;
		15'h0726: char_row_bitmap <= 16'b0000001100000000;
		15'h0727: char_row_bitmap <= 16'b0000001100000000;
		15'h0728: char_row_bitmap <= 16'b0000001100000000;
		15'h0729: char_row_bitmap <= 16'b0000001100000000;
		15'h072a: char_row_bitmap <= 16'b0000001100000000;
		15'h072b: char_row_bitmap <= 16'b0000001111110000;
		15'h072c: char_row_bitmap <= 16'b0000001111110000;
		15'h072d: char_row_bitmap <= 16'b0000000000000000;
		15'h072e: char_row_bitmap <= 16'b0000000000000000;
		15'h072f: char_row_bitmap <= 16'b0000000000000000;
		15'h0730: char_row_bitmap <= 16'b1100000000000000;
		15'h0731: char_row_bitmap <= 16'b1110000000000000;
		15'h0732: char_row_bitmap <= 16'b0110000000000000;
		15'h0733: char_row_bitmap <= 16'b0011000000000000;
		15'h0734: char_row_bitmap <= 16'b0011100000000000;
		15'h0735: char_row_bitmap <= 16'b0001110000000000;
		15'h0736: char_row_bitmap <= 16'b0000111000000000;
		15'h0737: char_row_bitmap <= 16'b0000011000000000;
		15'h0738: char_row_bitmap <= 16'b0000011100000000;
		15'h0739: char_row_bitmap <= 16'b0000001110000000;
		15'h073a: char_row_bitmap <= 16'b0000000111000000;
		15'h073b: char_row_bitmap <= 16'b0000000011100000;
		15'h073c: char_row_bitmap <= 16'b0000000001100000;
		15'h073d: char_row_bitmap <= 16'b0000000001110000;
		15'h073e: char_row_bitmap <= 16'b0000000000111000;
		15'h073f: char_row_bitmap <= 16'b0000000000011100;
		15'h0740: char_row_bitmap <= 16'b0000000000001110;
		15'h0741: char_row_bitmap <= 16'b0000000000000110;
		15'h0742: char_row_bitmap <= 16'b0000000000000111;
		15'h0743: char_row_bitmap <= 16'b0000000000000011;
		15'h0744: char_row_bitmap <= 16'b0000000000000000;
		15'h0745: char_row_bitmap <= 16'b0000000000000000;
		15'h0746: char_row_bitmap <= 16'b0000111111000000;
		15'h0747: char_row_bitmap <= 16'b0000111111000000;
		15'h0748: char_row_bitmap <= 16'b0000000011000000;
		15'h0749: char_row_bitmap <= 16'b0000000011000000;
		15'h074a: char_row_bitmap <= 16'b0000000011000000;
		15'h074b: char_row_bitmap <= 16'b0000000011000000;
		15'h074c: char_row_bitmap <= 16'b0000000011000000;
		15'h074d: char_row_bitmap <= 16'b0000000011000000;
		15'h074e: char_row_bitmap <= 16'b0000000011000000;
		15'h074f: char_row_bitmap <= 16'b0000000011000000;
		15'h0750: char_row_bitmap <= 16'b0000000011000000;
		15'h0751: char_row_bitmap <= 16'b0000000011000000;
		15'h0752: char_row_bitmap <= 16'b0000000011000000;
		15'h0753: char_row_bitmap <= 16'b0000111111000000;
		15'h0754: char_row_bitmap <= 16'b0000111111000000;
		15'h0755: char_row_bitmap <= 16'b0000000000000000;
		15'h0756: char_row_bitmap <= 16'b0000000000000000;
		15'h0757: char_row_bitmap <= 16'b0000000000000000;
		15'h0758: char_row_bitmap <= 16'b0000000000000000;
		15'h0759: char_row_bitmap <= 16'b0000000000000000;
		15'h075a: char_row_bitmap <= 16'b0000001100000000;
		15'h075b: char_row_bitmap <= 16'b0000011110000000;
		15'h075c: char_row_bitmap <= 16'b0000111111000000;
		15'h075d: char_row_bitmap <= 16'b0001110011100000;
		15'h075e: char_row_bitmap <= 16'b0011100001110000;
		15'h075f: char_row_bitmap <= 16'b0011000000110000;
		15'h0760: char_row_bitmap <= 16'b0000000000000000;
		15'h0761: char_row_bitmap <= 16'b0000000000000000;
		15'h0762: char_row_bitmap <= 16'b0000000000000000;
		15'h0763: char_row_bitmap <= 16'b0000000000000000;
		15'h0764: char_row_bitmap <= 16'b0000000000000000;
		15'h0765: char_row_bitmap <= 16'b0000000000000000;
		15'h0766: char_row_bitmap <= 16'b0000000000000000;
		15'h0767: char_row_bitmap <= 16'b0000000000000000;
		15'h0768: char_row_bitmap <= 16'b0000000000000000;
		15'h0769: char_row_bitmap <= 16'b0000000000000000;
		15'h076a: char_row_bitmap <= 16'b0000000000000000;
		15'h076b: char_row_bitmap <= 16'b0000000000000000;
		15'h076c: char_row_bitmap <= 16'b0000000000000000;
		15'h076d: char_row_bitmap <= 16'b0000000000000000;
		15'h076e: char_row_bitmap <= 16'b0000000000000000;
		15'h076f: char_row_bitmap <= 16'b0000000000000000;
		15'h0770: char_row_bitmap <= 16'b0000000000000000;
		15'h0771: char_row_bitmap <= 16'b0000000000000000;
		15'h0772: char_row_bitmap <= 16'b0000000000000000;
		15'h0773: char_row_bitmap <= 16'b0000000000000000;
		15'h0774: char_row_bitmap <= 16'b0000000000000000;
		15'h0775: char_row_bitmap <= 16'b0000000000000000;
		15'h0776: char_row_bitmap <= 16'b0000000000000000;
		15'h0777: char_row_bitmap <= 16'b0000000000000000;
		15'h0778: char_row_bitmap <= 16'b0000000000000000;
		15'h0779: char_row_bitmap <= 16'b0000000000000000;
		15'h077a: char_row_bitmap <= 16'b0000000000000000;
		15'h077b: char_row_bitmap <= 16'b0000000000000000;
		15'h077c: char_row_bitmap <= 16'b0011111111111100;
		15'h077d: char_row_bitmap <= 16'b0011111111111100;
		15'h077e: char_row_bitmap <= 16'b0000000000000000;
		15'h077f: char_row_bitmap <= 16'b0000000000000000;
		15'h0780: char_row_bitmap <= 16'b0000000000000000;
		15'h0781: char_row_bitmap <= 16'b0000000000000000;
		15'h0782: char_row_bitmap <= 16'b0000001100000000;
		15'h0783: char_row_bitmap <= 16'b0000001100000000;
		15'h0784: char_row_bitmap <= 16'b0000001100000000;
		15'h0785: char_row_bitmap <= 16'b0000001110000000;
		15'h0786: char_row_bitmap <= 16'b0000000111000000;
		15'h0787: char_row_bitmap <= 16'b0000000011000000;
		15'h0788: char_row_bitmap <= 16'b0000000000000000;
		15'h0789: char_row_bitmap <= 16'b0000000000000000;
		15'h078a: char_row_bitmap <= 16'b0000000000000000;
		15'h078b: char_row_bitmap <= 16'b0000000000000000;
		15'h078c: char_row_bitmap <= 16'b0000000000000000;
		15'h078d: char_row_bitmap <= 16'b0000000000000000;
		15'h078e: char_row_bitmap <= 16'b0000000000000000;
		15'h078f: char_row_bitmap <= 16'b0000000000000000;
		15'h0790: char_row_bitmap <= 16'b0000000000000000;
		15'h0791: char_row_bitmap <= 16'b0000000000000000;
		15'h0792: char_row_bitmap <= 16'b0000000000000000;
		15'h0793: char_row_bitmap <= 16'b0000000000000000;
		15'h0794: char_row_bitmap <= 16'b0000000000000000;
		15'h0795: char_row_bitmap <= 16'b0000000000000000;
		15'h0796: char_row_bitmap <= 16'b0000000000000000;
		15'h0797: char_row_bitmap <= 16'b0000000000000000;
		15'h0798: char_row_bitmap <= 16'b0000000000000000;
		15'h0799: char_row_bitmap <= 16'b0000000000000000;
		15'h079a: char_row_bitmap <= 16'b0000111100110000;
		15'h079b: char_row_bitmap <= 16'b0001111110110000;
		15'h079c: char_row_bitmap <= 16'b0011100111110000;
		15'h079d: char_row_bitmap <= 16'b0011000011110000;
		15'h079e: char_row_bitmap <= 16'b0011000001110000;
		15'h079f: char_row_bitmap <= 16'b0011000001110000;
		15'h07a0: char_row_bitmap <= 16'b0011000011110000;
		15'h07a1: char_row_bitmap <= 16'b0011100111110000;
		15'h07a2: char_row_bitmap <= 16'b0001111110110000;
		15'h07a3: char_row_bitmap <= 16'b0000111100110000;
		15'h07a4: char_row_bitmap <= 16'b0000000000000000;
		15'h07a5: char_row_bitmap <= 16'b0000000000000000;
		15'h07a6: char_row_bitmap <= 16'b0000000000000000;
		15'h07a7: char_row_bitmap <= 16'b0000000000000000;
		15'h07a8: char_row_bitmap <= 16'b0000000000000000;
		15'h07a9: char_row_bitmap <= 16'b0000000000000000;
		15'h07aa: char_row_bitmap <= 16'b0011000000000000;
		15'h07ab: char_row_bitmap <= 16'b0011000000000000;
		15'h07ac: char_row_bitmap <= 16'b0011000000000000;
		15'h07ad: char_row_bitmap <= 16'b0011000000000000;
		15'h07ae: char_row_bitmap <= 16'b0011111111000000;
		15'h07af: char_row_bitmap <= 16'b0011111111100000;
		15'h07b0: char_row_bitmap <= 16'b0011000001110000;
		15'h07b1: char_row_bitmap <= 16'b0011000000110000;
		15'h07b2: char_row_bitmap <= 16'b0011000000110000;
		15'h07b3: char_row_bitmap <= 16'b0011000000110000;
		15'h07b4: char_row_bitmap <= 16'b0011000000110000;
		15'h07b5: char_row_bitmap <= 16'b0011000001110000;
		15'h07b6: char_row_bitmap <= 16'b0011111111100000;
		15'h07b7: char_row_bitmap <= 16'b0011111111000000;
		15'h07b8: char_row_bitmap <= 16'b0000000000000000;
		15'h07b9: char_row_bitmap <= 16'b0000000000000000;
		15'h07ba: char_row_bitmap <= 16'b0000000000000000;
		15'h07bb: char_row_bitmap <= 16'b0000000000000000;
		15'h07bc: char_row_bitmap <= 16'b0000000000000000;
		15'h07bd: char_row_bitmap <= 16'b0000000000000000;
		15'h07be: char_row_bitmap <= 16'b0000000000000000;
		15'h07bf: char_row_bitmap <= 16'b0000000000000000;
		15'h07c0: char_row_bitmap <= 16'b0000000000000000;
		15'h07c1: char_row_bitmap <= 16'b0000000000000000;
		15'h07c2: char_row_bitmap <= 16'b0000111111000000;
		15'h07c3: char_row_bitmap <= 16'b0001111111000000;
		15'h07c4: char_row_bitmap <= 16'b0011100000000000;
		15'h07c5: char_row_bitmap <= 16'b0011000000000000;
		15'h07c6: char_row_bitmap <= 16'b0011000000000000;
		15'h07c7: char_row_bitmap <= 16'b0011000000000000;
		15'h07c8: char_row_bitmap <= 16'b0011000000000000;
		15'h07c9: char_row_bitmap <= 16'b0011100000000000;
		15'h07ca: char_row_bitmap <= 16'b0001111111000000;
		15'h07cb: char_row_bitmap <= 16'b0000111111000000;
		15'h07cc: char_row_bitmap <= 16'b0000000000000000;
		15'h07cd: char_row_bitmap <= 16'b0000000000000000;
		15'h07ce: char_row_bitmap <= 16'b0000000000000000;
		15'h07cf: char_row_bitmap <= 16'b0000000000000000;
		15'h07d0: char_row_bitmap <= 16'b0000000000000000;
		15'h07d1: char_row_bitmap <= 16'b0000000000000000;
		15'h07d2: char_row_bitmap <= 16'b0000000000110000;
		15'h07d3: char_row_bitmap <= 16'b0000000000110000;
		15'h07d4: char_row_bitmap <= 16'b0000000000110000;
		15'h07d5: char_row_bitmap <= 16'b0000000000110000;
		15'h07d6: char_row_bitmap <= 16'b0000111111110000;
		15'h07d7: char_row_bitmap <= 16'b0001111111110000;
		15'h07d8: char_row_bitmap <= 16'b0011100000110000;
		15'h07d9: char_row_bitmap <= 16'b0011000000110000;
		15'h07da: char_row_bitmap <= 16'b0011000000110000;
		15'h07db: char_row_bitmap <= 16'b0011000000110000;
		15'h07dc: char_row_bitmap <= 16'b0011000000110000;
		15'h07dd: char_row_bitmap <= 16'b0011100000110000;
		15'h07de: char_row_bitmap <= 16'b0001111111110000;
		15'h07df: char_row_bitmap <= 16'b0000111111110000;
		15'h07e0: char_row_bitmap <= 16'b0000000000000000;
		15'h07e1: char_row_bitmap <= 16'b0000000000000000;
		15'h07e2: char_row_bitmap <= 16'b0000000000000000;
		15'h07e3: char_row_bitmap <= 16'b0000000000000000;
		15'h07e4: char_row_bitmap <= 16'b0000000000000000;
		15'h07e5: char_row_bitmap <= 16'b0000000000000000;
		15'h07e6: char_row_bitmap <= 16'b0000000000000000;
		15'h07e7: char_row_bitmap <= 16'b0000000000000000;
		15'h07e8: char_row_bitmap <= 16'b0000000000000000;
		15'h07e9: char_row_bitmap <= 16'b0000000000000000;
		15'h07ea: char_row_bitmap <= 16'b0000111111000000;
		15'h07eb: char_row_bitmap <= 16'b0001111111100000;
		15'h07ec: char_row_bitmap <= 16'b0011100001110000;
		15'h07ed: char_row_bitmap <= 16'b0011000000110000;
		15'h07ee: char_row_bitmap <= 16'b0011111111110000;
		15'h07ef: char_row_bitmap <= 16'b0011111111110000;
		15'h07f0: char_row_bitmap <= 16'b0011000000000000;
		15'h07f1: char_row_bitmap <= 16'b0011100000000000;
		15'h07f2: char_row_bitmap <= 16'b0001111111100000;
		15'h07f3: char_row_bitmap <= 16'b0000111111100000;
		15'h07f4: char_row_bitmap <= 16'b0000000000000000;
		15'h07f5: char_row_bitmap <= 16'b0000000000000000;
		15'h07f6: char_row_bitmap <= 16'b0000000000000000;
		15'h07f7: char_row_bitmap <= 16'b0000000000000000;
		15'h07f8: char_row_bitmap <= 16'b0000000000000000;
		15'h07f9: char_row_bitmap <= 16'b0000000000000000;
		15'h07fa: char_row_bitmap <= 16'b0000001111000000;
		15'h07fb: char_row_bitmap <= 16'b0000011111100000;
		15'h07fc: char_row_bitmap <= 16'b0000111001110000;
		15'h07fd: char_row_bitmap <= 16'b0000110000110000;
		15'h07fe: char_row_bitmap <= 16'b0000110000000000;
		15'h07ff: char_row_bitmap <= 16'b0000110000000000;
		15'h0800: char_row_bitmap <= 16'b0011111100000000;
		15'h0801: char_row_bitmap <= 16'b0011111100000000;
		15'h0802: char_row_bitmap <= 16'b0000110000000000;
		15'h0803: char_row_bitmap <= 16'b0000110000000000;
		15'h0804: char_row_bitmap <= 16'b0000110000000000;
		15'h0805: char_row_bitmap <= 16'b0000110000000000;
		15'h0806: char_row_bitmap <= 16'b0000110000000000;
		15'h0807: char_row_bitmap <= 16'b0000110000000000;
		15'h0808: char_row_bitmap <= 16'b0000000000000000;
		15'h0809: char_row_bitmap <= 16'b0000000000000000;
		15'h080a: char_row_bitmap <= 16'b0000000000000000;
		15'h080b: char_row_bitmap <= 16'b0000000000000000;
		15'h080c: char_row_bitmap <= 16'b0000000000000000;
		15'h080d: char_row_bitmap <= 16'b0000000000000000;
		15'h080e: char_row_bitmap <= 16'b0000000000000000;
		15'h080f: char_row_bitmap <= 16'b0000000000000000;
		15'h0810: char_row_bitmap <= 16'b0000000000000000;
		15'h0811: char_row_bitmap <= 16'b0000000000000000;
		15'h0812: char_row_bitmap <= 16'b0000111111110000;
		15'h0813: char_row_bitmap <= 16'b0001111111110000;
		15'h0814: char_row_bitmap <= 16'b0011100000110000;
		15'h0815: char_row_bitmap <= 16'b0011000000110000;
		15'h0816: char_row_bitmap <= 16'b0011000000110000;
		15'h0817: char_row_bitmap <= 16'b0011100000110000;
		15'h0818: char_row_bitmap <= 16'b0001111111110000;
		15'h0819: char_row_bitmap <= 16'b0000111111110000;
		15'h081a: char_row_bitmap <= 16'b0000000000110000;
		15'h081b: char_row_bitmap <= 16'b0000000000110000;
		15'h081c: char_row_bitmap <= 16'b0001100000110000;
		15'h081d: char_row_bitmap <= 16'b0001110001110000;
		15'h081e: char_row_bitmap <= 16'b0000111111100000;
		15'h081f: char_row_bitmap <= 16'b0000011111000000;
		15'h0820: char_row_bitmap <= 16'b0000000000000000;
		15'h0821: char_row_bitmap <= 16'b0000000000000000;
		15'h0822: char_row_bitmap <= 16'b0011000000000000;
		15'h0823: char_row_bitmap <= 16'b0011000000000000;
		15'h0824: char_row_bitmap <= 16'b0011000000000000;
		15'h0825: char_row_bitmap <= 16'b0011000000000000;
		15'h0826: char_row_bitmap <= 16'b0011001111000000;
		15'h0827: char_row_bitmap <= 16'b0011011111100000;
		15'h0828: char_row_bitmap <= 16'b0011111001110000;
		15'h0829: char_row_bitmap <= 16'b0011110000110000;
		15'h082a: char_row_bitmap <= 16'b0011100000110000;
		15'h082b: char_row_bitmap <= 16'b0011000000110000;
		15'h082c: char_row_bitmap <= 16'b0011000000110000;
		15'h082d: char_row_bitmap <= 16'b0011000000110000;
		15'h082e: char_row_bitmap <= 16'b0011000000110000;
		15'h082f: char_row_bitmap <= 16'b0011000000110000;
		15'h0830: char_row_bitmap <= 16'b0000000000000000;
		15'h0831: char_row_bitmap <= 16'b0000000000000000;
		15'h0832: char_row_bitmap <= 16'b0000000000000000;
		15'h0833: char_row_bitmap <= 16'b0000000000000000;
		15'h0834: char_row_bitmap <= 16'b0000000000000000;
		15'h0835: char_row_bitmap <= 16'b0000000000000000;
		15'h0836: char_row_bitmap <= 16'b0000001100000000;
		15'h0837: char_row_bitmap <= 16'b0000001100000000;
		15'h0838: char_row_bitmap <= 16'b0000000000000000;
		15'h0839: char_row_bitmap <= 16'b0000000000000000;
		15'h083a: char_row_bitmap <= 16'b0000111100000000;
		15'h083b: char_row_bitmap <= 16'b0000111100000000;
		15'h083c: char_row_bitmap <= 16'b0000001100000000;
		15'h083d: char_row_bitmap <= 16'b0000001100000000;
		15'h083e: char_row_bitmap <= 16'b0000001100000000;
		15'h083f: char_row_bitmap <= 16'b0000001100000000;
		15'h0840: char_row_bitmap <= 16'b0000001100000000;
		15'h0841: char_row_bitmap <= 16'b0000001100000000;
		15'h0842: char_row_bitmap <= 16'b0000111111000000;
		15'h0843: char_row_bitmap <= 16'b0000111111000000;
		15'h0844: char_row_bitmap <= 16'b0000000000000000;
		15'h0845: char_row_bitmap <= 16'b0000000000000000;
		15'h0846: char_row_bitmap <= 16'b0000000000000000;
		15'h0847: char_row_bitmap <= 16'b0000000000000000;
		15'h0848: char_row_bitmap <= 16'b0000000000000000;
		15'h0849: char_row_bitmap <= 16'b0000000000000000;
		15'h084a: char_row_bitmap <= 16'b0000000011000000;
		15'h084b: char_row_bitmap <= 16'b0000000011000000;
		15'h084c: char_row_bitmap <= 16'b0000000000000000;
		15'h084d: char_row_bitmap <= 16'b0000000000000000;
		15'h084e: char_row_bitmap <= 16'b0000001111000000;
		15'h084f: char_row_bitmap <= 16'b0000001111000000;
		15'h0850: char_row_bitmap <= 16'b0000000011000000;
		15'h0851: char_row_bitmap <= 16'b0000000011000000;
		15'h0852: char_row_bitmap <= 16'b0000000011000000;
		15'h0853: char_row_bitmap <= 16'b0000000011000000;
		15'h0854: char_row_bitmap <= 16'b0000000011000000;
		15'h0855: char_row_bitmap <= 16'b0000000011000000;
		15'h0856: char_row_bitmap <= 16'b0000000011000000;
		15'h0857: char_row_bitmap <= 16'b0000000011000000;
		15'h0858: char_row_bitmap <= 16'b0011000011000000;
		15'h0859: char_row_bitmap <= 16'b0011100111000000;
		15'h085a: char_row_bitmap <= 16'b0001111110000000;
		15'h085b: char_row_bitmap <= 16'b0000111100000000;
		15'h085c: char_row_bitmap <= 16'b0000000000000000;
		15'h085d: char_row_bitmap <= 16'b0000000000000000;
		15'h085e: char_row_bitmap <= 16'b0000110000000000;
		15'h085f: char_row_bitmap <= 16'b0000110000000000;
		15'h0860: char_row_bitmap <= 16'b0000110000000000;
		15'h0861: char_row_bitmap <= 16'b0000110000000000;
		15'h0862: char_row_bitmap <= 16'b0000110000110000;
		15'h0863: char_row_bitmap <= 16'b0000110001110000;
		15'h0864: char_row_bitmap <= 16'b0000110011100000;
		15'h0865: char_row_bitmap <= 16'b0000110111000000;
		15'h0866: char_row_bitmap <= 16'b0000111110000000;
		15'h0867: char_row_bitmap <= 16'b0000111110000000;
		15'h0868: char_row_bitmap <= 16'b0000110111000000;
		15'h0869: char_row_bitmap <= 16'b0000110011100000;
		15'h086a: char_row_bitmap <= 16'b0000110001110000;
		15'h086b: char_row_bitmap <= 16'b0000110000110000;
		15'h086c: char_row_bitmap <= 16'b0000000000000000;
		15'h086d: char_row_bitmap <= 16'b0000000000000000;
		15'h086e: char_row_bitmap <= 16'b0000000000000000;
		15'h086f: char_row_bitmap <= 16'b0000000000000000;
		15'h0870: char_row_bitmap <= 16'b0000000000000000;
		15'h0871: char_row_bitmap <= 16'b0000000000000000;
		15'h0872: char_row_bitmap <= 16'b0000111100000000;
		15'h0873: char_row_bitmap <= 16'b0000111100000000;
		15'h0874: char_row_bitmap <= 16'b0000001100000000;
		15'h0875: char_row_bitmap <= 16'b0000001100000000;
		15'h0876: char_row_bitmap <= 16'b0000001100000000;
		15'h0877: char_row_bitmap <= 16'b0000001100000000;
		15'h0878: char_row_bitmap <= 16'b0000001100000000;
		15'h0879: char_row_bitmap <= 16'b0000001100000000;
		15'h087a: char_row_bitmap <= 16'b0000001100000000;
		15'h087b: char_row_bitmap <= 16'b0000001100000000;
		15'h087c: char_row_bitmap <= 16'b0000001100000000;
		15'h087d: char_row_bitmap <= 16'b0000001100000000;
		15'h087e: char_row_bitmap <= 16'b0000111111000000;
		15'h087f: char_row_bitmap <= 16'b0000111111000000;
		15'h0880: char_row_bitmap <= 16'b0000000000000000;
		15'h0881: char_row_bitmap <= 16'b0000000000000000;
		15'h0882: char_row_bitmap <= 16'b0000000000000000;
		15'h0883: char_row_bitmap <= 16'b0000000000000000;
		15'h0884: char_row_bitmap <= 16'b0000000000000000;
		15'h0885: char_row_bitmap <= 16'b0000000000000000;
		15'h0886: char_row_bitmap <= 16'b0000000000000000;
		15'h0887: char_row_bitmap <= 16'b0000000000000000;
		15'h0888: char_row_bitmap <= 16'b0000000000000000;
		15'h0889: char_row_bitmap <= 16'b0000000000000000;
		15'h088a: char_row_bitmap <= 16'b0011110011000000;
		15'h088b: char_row_bitmap <= 16'b0011111111100000;
		15'h088c: char_row_bitmap <= 16'b0011111111110000;
		15'h088d: char_row_bitmap <= 16'b0011001100110000;
		15'h088e: char_row_bitmap <= 16'b0011001100110000;
		15'h088f: char_row_bitmap <= 16'b0011001100110000;
		15'h0890: char_row_bitmap <= 16'b0011001100110000;
		15'h0891: char_row_bitmap <= 16'b0011001100110000;
		15'h0892: char_row_bitmap <= 16'b0011001100110000;
		15'h0893: char_row_bitmap <= 16'b0011001100110000;
		15'h0894: char_row_bitmap <= 16'b0000000000000000;
		15'h0895: char_row_bitmap <= 16'b0000000000000000;
		15'h0896: char_row_bitmap <= 16'b0000000000000000;
		15'h0897: char_row_bitmap <= 16'b0000000000000000;
		15'h0898: char_row_bitmap <= 16'b0000000000000000;
		15'h0899: char_row_bitmap <= 16'b0000000000000000;
		15'h089a: char_row_bitmap <= 16'b0000000000000000;
		15'h089b: char_row_bitmap <= 16'b0000000000000000;
		15'h089c: char_row_bitmap <= 16'b0000000000000000;
		15'h089d: char_row_bitmap <= 16'b0000000000000000;
		15'h089e: char_row_bitmap <= 16'b0011001111000000;
		15'h089f: char_row_bitmap <= 16'b0011011111100000;
		15'h08a0: char_row_bitmap <= 16'b0011111001110000;
		15'h08a1: char_row_bitmap <= 16'b0011110000110000;
		15'h08a2: char_row_bitmap <= 16'b0011100000110000;
		15'h08a3: char_row_bitmap <= 16'b0011000000110000;
		15'h08a4: char_row_bitmap <= 16'b0011000000110000;
		15'h08a5: char_row_bitmap <= 16'b0011000000110000;
		15'h08a6: char_row_bitmap <= 16'b0011000000110000;
		15'h08a7: char_row_bitmap <= 16'b0011000000110000;
		15'h08a8: char_row_bitmap <= 16'b0000000000000000;
		15'h08a9: char_row_bitmap <= 16'b0000000000000000;
		15'h08aa: char_row_bitmap <= 16'b0000000000000000;
		15'h08ab: char_row_bitmap <= 16'b0000000000000000;
		15'h08ac: char_row_bitmap <= 16'b0000000000000000;
		15'h08ad: char_row_bitmap <= 16'b0000000000000000;
		15'h08ae: char_row_bitmap <= 16'b0000000000000000;
		15'h08af: char_row_bitmap <= 16'b0000000000000000;
		15'h08b0: char_row_bitmap <= 16'b0000000000000000;
		15'h08b1: char_row_bitmap <= 16'b0000000000000000;
		15'h08b2: char_row_bitmap <= 16'b0000111111000000;
		15'h08b3: char_row_bitmap <= 16'b0001111111100000;
		15'h08b4: char_row_bitmap <= 16'b0011100001110000;
		15'h08b5: char_row_bitmap <= 16'b0011000000110000;
		15'h08b6: char_row_bitmap <= 16'b0011000000110000;
		15'h08b7: char_row_bitmap <= 16'b0011000000110000;
		15'h08b8: char_row_bitmap <= 16'b0011000000110000;
		15'h08b9: char_row_bitmap <= 16'b0011100001110000;
		15'h08ba: char_row_bitmap <= 16'b0001111111100000;
		15'h08bb: char_row_bitmap <= 16'b0000111111000000;
		15'h08bc: char_row_bitmap <= 16'b0000000000000000;
		15'h08bd: char_row_bitmap <= 16'b0000000000000000;
		15'h08be: char_row_bitmap <= 16'b0000000000000000;
		15'h08bf: char_row_bitmap <= 16'b0000000000000000;
		15'h08c0: char_row_bitmap <= 16'b0000000000000000;
		15'h08c1: char_row_bitmap <= 16'b0000000000000000;
		15'h08c2: char_row_bitmap <= 16'b0000000000000000;
		15'h08c3: char_row_bitmap <= 16'b0000000000000000;
		15'h08c4: char_row_bitmap <= 16'b0000000000000000;
		15'h08c5: char_row_bitmap <= 16'b0000000000000000;
		15'h08c6: char_row_bitmap <= 16'b0011111111000000;
		15'h08c7: char_row_bitmap <= 16'b0011111111100000;
		15'h08c8: char_row_bitmap <= 16'b0011000001110000;
		15'h08c9: char_row_bitmap <= 16'b0011000000110000;
		15'h08ca: char_row_bitmap <= 16'b0011000000110000;
		15'h08cb: char_row_bitmap <= 16'b0011000000110000;
		15'h08cc: char_row_bitmap <= 16'b0011000000110000;
		15'h08cd: char_row_bitmap <= 16'b0011000001110000;
		15'h08ce: char_row_bitmap <= 16'b0011111111100000;
		15'h08cf: char_row_bitmap <= 16'b0011111111000000;
		15'h08d0: char_row_bitmap <= 16'b0011000000000000;
		15'h08d1: char_row_bitmap <= 16'b0011000000000000;
		15'h08d2: char_row_bitmap <= 16'b0011000000000000;
		15'h08d3: char_row_bitmap <= 16'b0011000000000000;
		15'h08d4: char_row_bitmap <= 16'b0000000000000000;
		15'h08d5: char_row_bitmap <= 16'b0000000000000000;
		15'h08d6: char_row_bitmap <= 16'b0000000000000000;
		15'h08d7: char_row_bitmap <= 16'b0000000000000000;
		15'h08d8: char_row_bitmap <= 16'b0000000000000000;
		15'h08d9: char_row_bitmap <= 16'b0000000000000000;
		15'h08da: char_row_bitmap <= 16'b0000111111110000;
		15'h08db: char_row_bitmap <= 16'b0001111111110000;
		15'h08dc: char_row_bitmap <= 16'b0011100000110000;
		15'h08dd: char_row_bitmap <= 16'b0011000000110000;
		15'h08de: char_row_bitmap <= 16'b0011000000110000;
		15'h08df: char_row_bitmap <= 16'b0011000000110000;
		15'h08e0: char_row_bitmap <= 16'b0011000000110000;
		15'h08e1: char_row_bitmap <= 16'b0011100000110000;
		15'h08e2: char_row_bitmap <= 16'b0001111111110000;
		15'h08e3: char_row_bitmap <= 16'b0000111111110000;
		15'h08e4: char_row_bitmap <= 16'b0000000000110000;
		15'h08e5: char_row_bitmap <= 16'b0000000000110000;
		15'h08e6: char_row_bitmap <= 16'b0000000000110000;
		15'h08e7: char_row_bitmap <= 16'b0000000000110000;
		15'h08e8: char_row_bitmap <= 16'b0000000000000000;
		15'h08e9: char_row_bitmap <= 16'b0000000000000000;
		15'h08ea: char_row_bitmap <= 16'b0000000000000000;
		15'h08eb: char_row_bitmap <= 16'b0000000000000000;
		15'h08ec: char_row_bitmap <= 16'b0000000000000000;
		15'h08ed: char_row_bitmap <= 16'b0000000000000000;
		15'h08ee: char_row_bitmap <= 16'b0011001111000000;
		15'h08ef: char_row_bitmap <= 16'b0011011111100000;
		15'h08f0: char_row_bitmap <= 16'b0011111001110000;
		15'h08f1: char_row_bitmap <= 16'b0011110000110000;
		15'h08f2: char_row_bitmap <= 16'b0011100000000000;
		15'h08f3: char_row_bitmap <= 16'b0011000000000000;
		15'h08f4: char_row_bitmap <= 16'b0011000000000000;
		15'h08f5: char_row_bitmap <= 16'b0011000000000000;
		15'h08f6: char_row_bitmap <= 16'b0011000000000000;
		15'h08f7: char_row_bitmap <= 16'b0011000000000000;
		15'h08f8: char_row_bitmap <= 16'b0000000000000000;
		15'h08f9: char_row_bitmap <= 16'b0000000000000000;
		15'h08fa: char_row_bitmap <= 16'b0000000000000000;
		15'h08fb: char_row_bitmap <= 16'b0000000000000000;
		15'h08fc: char_row_bitmap <= 16'b0000000000000000;
		15'h08fd: char_row_bitmap <= 16'b0000000000000000;
		15'h08fe: char_row_bitmap <= 16'b0000000000000000;
		15'h08ff: char_row_bitmap <= 16'b0000000000000000;
		15'h0900: char_row_bitmap <= 16'b0000000000000000;
		15'h0901: char_row_bitmap <= 16'b0000000000000000;
		15'h0902: char_row_bitmap <= 16'b0000111111100000;
		15'h0903: char_row_bitmap <= 16'b0001111111100000;
		15'h0904: char_row_bitmap <= 16'b0011100000000000;
		15'h0905: char_row_bitmap <= 16'b0011100000000000;
		15'h0906: char_row_bitmap <= 16'b0001111111000000;
		15'h0907: char_row_bitmap <= 16'b0000111111100000;
		15'h0908: char_row_bitmap <= 16'b0000000001110000;
		15'h0909: char_row_bitmap <= 16'b0000000001110000;
		15'h090a: char_row_bitmap <= 16'b0011111111100000;
		15'h090b: char_row_bitmap <= 16'b0011111111000000;
		15'h090c: char_row_bitmap <= 16'b0000000000000000;
		15'h090d: char_row_bitmap <= 16'b0000000000000000;
		15'h090e: char_row_bitmap <= 16'b0000000000000000;
		15'h090f: char_row_bitmap <= 16'b0000000000000000;
		15'h0910: char_row_bitmap <= 16'b0000000000000000;
		15'h0911: char_row_bitmap <= 16'b0000000000000000;
		15'h0912: char_row_bitmap <= 16'b0000110000000000;
		15'h0913: char_row_bitmap <= 16'b0000110000000000;
		15'h0914: char_row_bitmap <= 16'b0000110000000000;
		15'h0915: char_row_bitmap <= 16'b0000110000000000;
		15'h0916: char_row_bitmap <= 16'b0000111111000000;
		15'h0917: char_row_bitmap <= 16'b0000111111000000;
		15'h0918: char_row_bitmap <= 16'b0000110000000000;
		15'h0919: char_row_bitmap <= 16'b0000110000000000;
		15'h091a: char_row_bitmap <= 16'b0000110000000000;
		15'h091b: char_row_bitmap <= 16'b0000110000000000;
		15'h091c: char_row_bitmap <= 16'b0000110000000000;
		15'h091d: char_row_bitmap <= 16'b0000111000000000;
		15'h091e: char_row_bitmap <= 16'b0000011111000000;
		15'h091f: char_row_bitmap <= 16'b0000001111000000;
		15'h0920: char_row_bitmap <= 16'b0000000000000000;
		15'h0921: char_row_bitmap <= 16'b0000000000000000;
		15'h0922: char_row_bitmap <= 16'b0000000000000000;
		15'h0923: char_row_bitmap <= 16'b0000000000000000;
		15'h0924: char_row_bitmap <= 16'b0000000000000000;
		15'h0925: char_row_bitmap <= 16'b0000000000000000;
		15'h0926: char_row_bitmap <= 16'b0000000000000000;
		15'h0927: char_row_bitmap <= 16'b0000000000000000;
		15'h0928: char_row_bitmap <= 16'b0000000000000000;
		15'h0929: char_row_bitmap <= 16'b0000000000000000;
		15'h092a: char_row_bitmap <= 16'b0011000000110000;
		15'h092b: char_row_bitmap <= 16'b0011000000110000;
		15'h092c: char_row_bitmap <= 16'b0011000000110000;
		15'h092d: char_row_bitmap <= 16'b0011000000110000;
		15'h092e: char_row_bitmap <= 16'b0011000000110000;
		15'h092f: char_row_bitmap <= 16'b0011000001110000;
		15'h0930: char_row_bitmap <= 16'b0011000011110000;
		15'h0931: char_row_bitmap <= 16'b0011100111110000;
		15'h0932: char_row_bitmap <= 16'b0001111110110000;
		15'h0933: char_row_bitmap <= 16'b0000111100110000;
		15'h0934: char_row_bitmap <= 16'b0000000000000000;
		15'h0935: char_row_bitmap <= 16'b0000000000000000;
		15'h0936: char_row_bitmap <= 16'b0000000000000000;
		15'h0937: char_row_bitmap <= 16'b0000000000000000;
		15'h0938: char_row_bitmap <= 16'b0000000000000000;
		15'h0939: char_row_bitmap <= 16'b0000000000000000;
		15'h093a: char_row_bitmap <= 16'b0000000000000000;
		15'h093b: char_row_bitmap <= 16'b0000000000000000;
		15'h093c: char_row_bitmap <= 16'b0000000000000000;
		15'h093d: char_row_bitmap <= 16'b0000000000000000;
		15'h093e: char_row_bitmap <= 16'b0011000000110000;
		15'h093f: char_row_bitmap <= 16'b0011000000110000;
		15'h0940: char_row_bitmap <= 16'b0011100001110000;
		15'h0941: char_row_bitmap <= 16'b0001100001100000;
		15'h0942: char_row_bitmap <= 16'b0001110011100000;
		15'h0943: char_row_bitmap <= 16'b0000110011000000;
		15'h0944: char_row_bitmap <= 16'b0000110011000000;
		15'h0945: char_row_bitmap <= 16'b0000011110000000;
		15'h0946: char_row_bitmap <= 16'b0000011110000000;
		15'h0947: char_row_bitmap <= 16'b0000001100000000;
		15'h0948: char_row_bitmap <= 16'b0000000000000000;
		15'h0949: char_row_bitmap <= 16'b0000000000000000;
		15'h094a: char_row_bitmap <= 16'b0000000000000000;
		15'h094b: char_row_bitmap <= 16'b0000000000000000;
		15'h094c: char_row_bitmap <= 16'b0000000000000000;
		15'h094d: char_row_bitmap <= 16'b0000000000000000;
		15'h094e: char_row_bitmap <= 16'b0000000000000000;
		15'h094f: char_row_bitmap <= 16'b0000000000000000;
		15'h0950: char_row_bitmap <= 16'b0000000000000000;
		15'h0951: char_row_bitmap <= 16'b0000000000000000;
		15'h0952: char_row_bitmap <= 16'b0011000000110000;
		15'h0953: char_row_bitmap <= 16'b0011000000110000;
		15'h0954: char_row_bitmap <= 16'b0011000000110000;
		15'h0955: char_row_bitmap <= 16'b0011000000110000;
		15'h0956: char_row_bitmap <= 16'b0011001100110000;
		15'h0957: char_row_bitmap <= 16'b0011001100110000;
		15'h0958: char_row_bitmap <= 16'b0011001100110000;
		15'h0959: char_row_bitmap <= 16'b0011111111110000;
		15'h095a: char_row_bitmap <= 16'b0001111111100000;
		15'h095b: char_row_bitmap <= 16'b0000110011000000;
		15'h095c: char_row_bitmap <= 16'b0000000000000000;
		15'h095d: char_row_bitmap <= 16'b0000000000000000;
		15'h095e: char_row_bitmap <= 16'b0000000000000000;
		15'h095f: char_row_bitmap <= 16'b0000000000000000;
		15'h0960: char_row_bitmap <= 16'b0000000000000000;
		15'h0961: char_row_bitmap <= 16'b0000000000000000;
		15'h0962: char_row_bitmap <= 16'b0000000000000000;
		15'h0963: char_row_bitmap <= 16'b0000000000000000;
		15'h0964: char_row_bitmap <= 16'b0000000000000000;
		15'h0965: char_row_bitmap <= 16'b0000000000000000;
		15'h0966: char_row_bitmap <= 16'b0011000000110000;
		15'h0967: char_row_bitmap <= 16'b0011100001110000;
		15'h0968: char_row_bitmap <= 16'b0001110011100000;
		15'h0969: char_row_bitmap <= 16'b0000111111000000;
		15'h096a: char_row_bitmap <= 16'b0000011110000000;
		15'h096b: char_row_bitmap <= 16'b0000011110000000;
		15'h096c: char_row_bitmap <= 16'b0000111111000000;
		15'h096d: char_row_bitmap <= 16'b0001110011100000;
		15'h096e: char_row_bitmap <= 16'b0011100001110000;
		15'h096f: char_row_bitmap <= 16'b0011000000110000;
		15'h0970: char_row_bitmap <= 16'b0000000000000000;
		15'h0971: char_row_bitmap <= 16'b0000000000000000;
		15'h0972: char_row_bitmap <= 16'b0000000000000000;
		15'h0973: char_row_bitmap <= 16'b0000000000000000;
		15'h0974: char_row_bitmap <= 16'b0000000000000000;
		15'h0975: char_row_bitmap <= 16'b0000000000000000;
		15'h0976: char_row_bitmap <= 16'b0000000000000000;
		15'h0977: char_row_bitmap <= 16'b0000000000000000;
		15'h0978: char_row_bitmap <= 16'b0000000000000000;
		15'h0979: char_row_bitmap <= 16'b0000000000000000;
		15'h097a: char_row_bitmap <= 16'b0011000000110000;
		15'h097b: char_row_bitmap <= 16'b0011000000110000;
		15'h097c: char_row_bitmap <= 16'b0011000000110000;
		15'h097d: char_row_bitmap <= 16'b0011000001110000;
		15'h097e: char_row_bitmap <= 16'b0011000011110000;
		15'h097f: char_row_bitmap <= 16'b0011100111110000;
		15'h0980: char_row_bitmap <= 16'b0001111110110000;
		15'h0981: char_row_bitmap <= 16'b0000111100110000;
		15'h0982: char_row_bitmap <= 16'b0000000000110000;
		15'h0983: char_row_bitmap <= 16'b0000000000110000;
		15'h0984: char_row_bitmap <= 16'b0011000000110000;
		15'h0985: char_row_bitmap <= 16'b0011100001110000;
		15'h0986: char_row_bitmap <= 16'b0001111111100000;
		15'h0987: char_row_bitmap <= 16'b0000111111000000;
		15'h0988: char_row_bitmap <= 16'b0000000000000000;
		15'h0989: char_row_bitmap <= 16'b0000000000000000;
		15'h098a: char_row_bitmap <= 16'b0000000000000000;
		15'h098b: char_row_bitmap <= 16'b0000000000000000;
		15'h098c: char_row_bitmap <= 16'b0000000000000000;
		15'h098d: char_row_bitmap <= 16'b0000000000000000;
		15'h098e: char_row_bitmap <= 16'b0011111111110000;
		15'h098f: char_row_bitmap <= 16'b0011111111110000;
		15'h0990: char_row_bitmap <= 16'b0000000011100000;
		15'h0991: char_row_bitmap <= 16'b0000000111000000;
		15'h0992: char_row_bitmap <= 16'b0000001110000000;
		15'h0993: char_row_bitmap <= 16'b0000011100000000;
		15'h0994: char_row_bitmap <= 16'b0000111000000000;
		15'h0995: char_row_bitmap <= 16'b0001110000000000;
		15'h0996: char_row_bitmap <= 16'b0011111111110000;
		15'h0997: char_row_bitmap <= 16'b0011111111110000;
		15'h0998: char_row_bitmap <= 16'b0000000000000000;
		15'h0999: char_row_bitmap <= 16'b0000000000000000;
		15'h099a: char_row_bitmap <= 16'b0000000000000000;
		15'h099b: char_row_bitmap <= 16'b0000000000000000;
		15'h099c: char_row_bitmap <= 16'b0000000000000000;
		15'h099d: char_row_bitmap <= 16'b0000000000000000;
		15'h099e: char_row_bitmap <= 16'b0000000011110000;
		15'h099f: char_row_bitmap <= 16'b0000000111110000;
		15'h09a0: char_row_bitmap <= 16'b0000001110000000;
		15'h09a1: char_row_bitmap <= 16'b0000001100000000;
		15'h09a2: char_row_bitmap <= 16'b0000001100000000;
		15'h09a3: char_row_bitmap <= 16'b0000011100000000;
		15'h09a4: char_row_bitmap <= 16'b0000111000000000;
		15'h09a5: char_row_bitmap <= 16'b0001110000000000;
		15'h09a6: char_row_bitmap <= 16'b0000111000000000;
		15'h09a7: char_row_bitmap <= 16'b0000011100000000;
		15'h09a8: char_row_bitmap <= 16'b0000001100000000;
		15'h09a9: char_row_bitmap <= 16'b0000001100000000;
		15'h09aa: char_row_bitmap <= 16'b0000001110000000;
		15'h09ab: char_row_bitmap <= 16'b0000000111110000;
		15'h09ac: char_row_bitmap <= 16'b0000000011110000;
		15'h09ad: char_row_bitmap <= 16'b0000000000000000;
		15'h09ae: char_row_bitmap <= 16'b0000000000000000;
		15'h09af: char_row_bitmap <= 16'b0000000000000000;
		15'h09b0: char_row_bitmap <= 16'b0000000000000000;
		15'h09b1: char_row_bitmap <= 16'b0000000000000000;
		15'h09b2: char_row_bitmap <= 16'b0000001100000000;
		15'h09b3: char_row_bitmap <= 16'b0000001100000000;
		15'h09b4: char_row_bitmap <= 16'b0000001100000000;
		15'h09b5: char_row_bitmap <= 16'b0000001100000000;
		15'h09b6: char_row_bitmap <= 16'b0000001100000000;
		15'h09b7: char_row_bitmap <= 16'b0000001100000000;
		15'h09b8: char_row_bitmap <= 16'b0000001100000000;
		15'h09b9: char_row_bitmap <= 16'b0000000000000000;
		15'h09ba: char_row_bitmap <= 16'b0000000000000000;
		15'h09bb: char_row_bitmap <= 16'b0000001100000000;
		15'h09bc: char_row_bitmap <= 16'b0000001100000000;
		15'h09bd: char_row_bitmap <= 16'b0000001100000000;
		15'h09be: char_row_bitmap <= 16'b0000001100000000;
		15'h09bf: char_row_bitmap <= 16'b0000001100000000;
		15'h09c0: char_row_bitmap <= 16'b0000001100000000;
		15'h09c1: char_row_bitmap <= 16'b0000001100000000;
		15'h09c2: char_row_bitmap <= 16'b0000000000000000;
		15'h09c3: char_row_bitmap <= 16'b0000000000000000;
		15'h09c4: char_row_bitmap <= 16'b0000000000000000;
		15'h09c5: char_row_bitmap <= 16'b0000000000000000;
		15'h09c6: char_row_bitmap <= 16'b0000111100000000;
		15'h09c7: char_row_bitmap <= 16'b0000111110000000;
		15'h09c8: char_row_bitmap <= 16'b0000000111000000;
		15'h09c9: char_row_bitmap <= 16'b0000000011000000;
		15'h09ca: char_row_bitmap <= 16'b0000000011000000;
		15'h09cb: char_row_bitmap <= 16'b0000000011100000;
		15'h09cc: char_row_bitmap <= 16'b0000000001110000;
		15'h09cd: char_row_bitmap <= 16'b0000000000111000;
		15'h09ce: char_row_bitmap <= 16'b0000000001110000;
		15'h09cf: char_row_bitmap <= 16'b0000000011100000;
		15'h09d0: char_row_bitmap <= 16'b0000000011000000;
		15'h09d1: char_row_bitmap <= 16'b0000000011000000;
		15'h09d2: char_row_bitmap <= 16'b0000000111000000;
		15'h09d3: char_row_bitmap <= 16'b0000111110000000;
		15'h09d4: char_row_bitmap <= 16'b0000111100000000;
		15'h09d5: char_row_bitmap <= 16'b0000000000000000;
		15'h09d6: char_row_bitmap <= 16'b0000000000000000;
		15'h09d7: char_row_bitmap <= 16'b0000000000000000;
		15'h09d8: char_row_bitmap <= 16'b0000000000000000;
		15'h09d9: char_row_bitmap <= 16'b0000000000000000;
		15'h09da: char_row_bitmap <= 16'b0000000000000000;
		15'h09db: char_row_bitmap <= 16'b0000000000000000;
		15'h09dc: char_row_bitmap <= 16'b0000000000000000;
		15'h09dd: char_row_bitmap <= 16'b0000000000000000;
		15'h09de: char_row_bitmap <= 16'b0000000000000000;
		15'h09df: char_row_bitmap <= 16'b0000000000000000;
		15'h09e0: char_row_bitmap <= 16'b0000111100001100;
		15'h09e1: char_row_bitmap <= 16'b0001111110011100;
		15'h09e2: char_row_bitmap <= 16'b0011100111111000;
		15'h09e3: char_row_bitmap <= 16'b0011000011110000;
		15'h09e4: char_row_bitmap <= 16'b0000000000000000;
		15'h09e5: char_row_bitmap <= 16'b0000000000000000;
		15'h09e6: char_row_bitmap <= 16'b0000000000000000;
		15'h09e7: char_row_bitmap <= 16'b0000000000000000;
		15'h09e8: char_row_bitmap <= 16'b0000000000000000;
		15'h09e9: char_row_bitmap <= 16'b0000000000000000;
		15'h09ea: char_row_bitmap <= 16'b0000000000000000;
		15'h09eb: char_row_bitmap <= 16'b0000000000000000;
		15'h09ec: char_row_bitmap <= 16'b0000000000000000;
		15'h09ed: char_row_bitmap <= 16'b0000000000000000;
		15'h09ee: char_row_bitmap <= 16'b0111111011000110;
		15'h09ef: char_row_bitmap <= 16'b0111111011101110;
		15'h09f0: char_row_bitmap <= 16'b0001100011111110;
		15'h09f1: char_row_bitmap <= 16'b0001100011010110;
		15'h09f2: char_row_bitmap <= 16'b0001100011000110;
		15'h09f3: char_row_bitmap <= 16'b0001100011000110;
		15'h09f4: char_row_bitmap <= 16'b0001100011000110;
		15'h09f5: char_row_bitmap <= 16'b0000000000000000;
		15'h09f6: char_row_bitmap <= 16'b0000000000000000;
		15'h09f7: char_row_bitmap <= 16'b0000000000000000;
		15'h09f8: char_row_bitmap <= 16'b0000000000000000;
		15'h09f9: char_row_bitmap <= 16'b0000000000000000;
		15'h09fa: char_row_bitmap <= 16'b0000000000000000;
		15'h09fb: char_row_bitmap <= 16'b0000000000000000;
		15'h09fc: char_row_bitmap <= 16'b0000000000000000;
		15'h09fd: char_row_bitmap <= 16'b0000000000000000;
		15'h09fe: char_row_bitmap <= 16'b0000000000000000;
		15'h09ff: char_row_bitmap <= 16'b0000000000000000;
		15'h0a00: char_row_bitmap <= 16'b0000000000000000;
		15'h0a01: char_row_bitmap <= 16'b0000000000000000;
		15'h0a02: char_row_bitmap <= 16'b0100100000000000;
		15'h0a03: char_row_bitmap <= 16'b0110100000000000;
		15'h0a04: char_row_bitmap <= 16'b0101100000000000;
		15'h0a05: char_row_bitmap <= 16'b0100100000000000;
		15'h0a06: char_row_bitmap <= 16'b0100100000000000;
		15'h0a07: char_row_bitmap <= 16'b0000000000000000;
		15'h0a08: char_row_bitmap <= 16'b0000001001000000;
		15'h0a09: char_row_bitmap <= 16'b0000001001000000;
		15'h0a0a: char_row_bitmap <= 16'b0000001001000000;
		15'h0a0b: char_row_bitmap <= 16'b0000001001000000;
		15'h0a0c: char_row_bitmap <= 16'b0000000110000000;
		15'h0a0d: char_row_bitmap <= 16'b0000000000000000;
		15'h0a0e: char_row_bitmap <= 16'b0000000000010000;
		15'h0a0f: char_row_bitmap <= 16'b0000000000010000;
		15'h0a10: char_row_bitmap <= 16'b0000000000010000;
		15'h0a11: char_row_bitmap <= 16'b0000000000010000;
		15'h0a12: char_row_bitmap <= 16'b0000000000011110;
		15'h0a13: char_row_bitmap <= 16'b0000000000000000;
		15'h0a14: char_row_bitmap <= 16'b0000000000000000;
		15'h0a15: char_row_bitmap <= 16'b0000000000000000;
		15'h0a16: char_row_bitmap <= 16'b0011100000000000;
		15'h0a17: char_row_bitmap <= 16'b0100000000000000;
		15'h0a18: char_row_bitmap <= 16'b0011000000000000;
		15'h0a19: char_row_bitmap <= 16'b0000100000000000;
		15'h0a1a: char_row_bitmap <= 16'b0111000000000000;
		15'h0a1b: char_row_bitmap <= 16'b0000000000000000;
		15'h0a1c: char_row_bitmap <= 16'b0000000110000000;
		15'h0a1d: char_row_bitmap <= 16'b0000001001000000;
		15'h0a1e: char_row_bitmap <= 16'b0000001001000000;
		15'h0a1f: char_row_bitmap <= 16'b0000001001000000;
		15'h0a20: char_row_bitmap <= 16'b0000000110000000;
		15'h0a21: char_row_bitmap <= 16'b0000000000000000;
		15'h0a22: char_row_bitmap <= 16'b0000000000010010;
		15'h0a23: char_row_bitmap <= 16'b0000000000010010;
		15'h0a24: char_row_bitmap <= 16'b0000000000011110;
		15'h0a25: char_row_bitmap <= 16'b0000000000010010;
		15'h0a26: char_row_bitmap <= 16'b0000000000010010;
		15'h0a27: char_row_bitmap <= 16'b0000000000000000;
		15'h0a28: char_row_bitmap <= 16'b0000000000000000;
		15'h0a29: char_row_bitmap <= 16'b0000000000000000;
		15'h0a2a: char_row_bitmap <= 16'b0011100000000000;
		15'h0a2b: char_row_bitmap <= 16'b0100000000000000;
		15'h0a2c: char_row_bitmap <= 16'b0011000000000000;
		15'h0a2d: char_row_bitmap <= 16'b0000100000000000;
		15'h0a2e: char_row_bitmap <= 16'b0111000000000000;
		15'h0a2f: char_row_bitmap <= 16'b0000000000000000;
		15'h0a30: char_row_bitmap <= 16'b0000001110000000;
		15'h0a31: char_row_bitmap <= 16'b0000000100000000;
		15'h0a32: char_row_bitmap <= 16'b0000000100000000;
		15'h0a33: char_row_bitmap <= 16'b0000000100000000;
		15'h0a34: char_row_bitmap <= 16'b0000000100000000;
		15'h0a35: char_row_bitmap <= 16'b0000000000000000;
		15'h0a36: char_row_bitmap <= 16'b0000000000100100;
		15'h0a37: char_row_bitmap <= 16'b0000000000100100;
		15'h0a38: char_row_bitmap <= 16'b0000000000011000;
		15'h0a39: char_row_bitmap <= 16'b0000000000100100;
		15'h0a3a: char_row_bitmap <= 16'b0000000000100100;
		15'h0a3b: char_row_bitmap <= 16'b0000000000000000;
		15'h0a3c: char_row_bitmap <= 16'b0000000000000000;
		15'h0a3d: char_row_bitmap <= 16'b0000000000000000;
		15'h0a3e: char_row_bitmap <= 16'b0111100000000000;
		15'h0a3f: char_row_bitmap <= 16'b0100000000000000;
		15'h0a40: char_row_bitmap <= 16'b0110000000000000;
		15'h0a41: char_row_bitmap <= 16'b0100000000000000;
		15'h0a42: char_row_bitmap <= 16'b0111100000000000;
		15'h0a43: char_row_bitmap <= 16'b0000000000000000;
		15'h0a44: char_row_bitmap <= 16'b0000001110000000;
		15'h0a45: char_row_bitmap <= 16'b0000000100000000;
		15'h0a46: char_row_bitmap <= 16'b0000000100000000;
		15'h0a47: char_row_bitmap <= 16'b0000000100000000;
		15'h0a48: char_row_bitmap <= 16'b0000000100000000;
		15'h0a49: char_row_bitmap <= 16'b0000000000000000;
		15'h0a4a: char_row_bitmap <= 16'b0000000000100100;
		15'h0a4b: char_row_bitmap <= 16'b0000000000100100;
		15'h0a4c: char_row_bitmap <= 16'b0000000000011000;
		15'h0a4d: char_row_bitmap <= 16'b0000000000100100;
		15'h0a4e: char_row_bitmap <= 16'b0000000000100100;
		15'h0a4f: char_row_bitmap <= 16'b0000000000000000;
		15'h0a50: char_row_bitmap <= 16'b0000000000000000;
		15'h0a51: char_row_bitmap <= 16'b0000000000000000;
		15'h0a52: char_row_bitmap <= 16'b0111100000000000;
		15'h0a53: char_row_bitmap <= 16'b0100000000000000;
		15'h0a54: char_row_bitmap <= 16'b0110000000000000;
		15'h0a55: char_row_bitmap <= 16'b0100000000000000;
		15'h0a56: char_row_bitmap <= 16'b0111100000000000;
		15'h0a57: char_row_bitmap <= 16'b0000000000000000;
		15'h0a58: char_row_bitmap <= 16'b0000000110000000;
		15'h0a59: char_row_bitmap <= 16'b0000001001000000;
		15'h0a5a: char_row_bitmap <= 16'b0000001001000000;
		15'h0a5b: char_row_bitmap <= 16'b0000001001000000;
		15'h0a5c: char_row_bitmap <= 16'b0000000110000000;
		15'h0a5d: char_row_bitmap <= 16'b0000000000000000;
		15'h0a5e: char_row_bitmap <= 16'b0000000000111000;
		15'h0a5f: char_row_bitmap <= 16'b0000000000010000;
		15'h0a60: char_row_bitmap <= 16'b0000000000010000;
		15'h0a61: char_row_bitmap <= 16'b0000000000010000;
		15'h0a62: char_row_bitmap <= 16'b0000000000010000;
		15'h0a63: char_row_bitmap <= 16'b0000000000000000;
		15'h0a64: char_row_bitmap <= 16'b0000000000000000;
		15'h0a65: char_row_bitmap <= 16'b0000000000000000;
		15'h0a66: char_row_bitmap <= 16'b0111100000000000;
		15'h0a67: char_row_bitmap <= 16'b0100000000000000;
		15'h0a68: char_row_bitmap <= 16'b0110000000000000;
		15'h0a69: char_row_bitmap <= 16'b0100000000000000;
		15'h0a6a: char_row_bitmap <= 16'b0111100000000000;
		15'h0a6b: char_row_bitmap <= 16'b0000000000000000;
		15'h0a6c: char_row_bitmap <= 16'b0000001001000000;
		15'h0a6d: char_row_bitmap <= 16'b0000001101000000;
		15'h0a6e: char_row_bitmap <= 16'b0000001011000000;
		15'h0a6f: char_row_bitmap <= 16'b0000001001000000;
		15'h0a70: char_row_bitmap <= 16'b0000001001000000;
		15'h0a71: char_row_bitmap <= 16'b0000000000000000;
		15'h0a72: char_row_bitmap <= 16'b0000000000001100;
		15'h0a73: char_row_bitmap <= 16'b0000000000010010;
		15'h0a74: char_row_bitmap <= 16'b0000000000010010;
		15'h0a75: char_row_bitmap <= 16'b0000000000010100;
		15'h0a76: char_row_bitmap <= 16'b0000000000001010;
		15'h0a77: char_row_bitmap <= 16'b0000000000000000;
		15'h0a78: char_row_bitmap <= 16'b0000000000000000;
		15'h0a79: char_row_bitmap <= 16'b0000000000000000;
		15'h0a7a: char_row_bitmap <= 16'b0011000000000000;
		15'h0a7b: char_row_bitmap <= 16'b0100100000000000;
		15'h0a7c: char_row_bitmap <= 16'b0111100000000000;
		15'h0a7d: char_row_bitmap <= 16'b0100100000000000;
		15'h0a7e: char_row_bitmap <= 16'b0100100000000000;
		15'h0a7f: char_row_bitmap <= 16'b0000000000000000;
		15'h0a80: char_row_bitmap <= 16'b0000000111000000;
		15'h0a81: char_row_bitmap <= 16'b0000001000000000;
		15'h0a82: char_row_bitmap <= 16'b0000001000000000;
		15'h0a83: char_row_bitmap <= 16'b0000001000000000;
		15'h0a84: char_row_bitmap <= 16'b0000000111000000;
		15'h0a85: char_row_bitmap <= 16'b0000000000000000;
		15'h0a86: char_row_bitmap <= 16'b0000000000010010;
		15'h0a87: char_row_bitmap <= 16'b0000000000010100;
		15'h0a88: char_row_bitmap <= 16'b0000000000011000;
		15'h0a89: char_row_bitmap <= 16'b0000000000010100;
		15'h0a8a: char_row_bitmap <= 16'b0000000000010010;
		15'h0a8b: char_row_bitmap <= 16'b0000000000000000;
		15'h0a8c: char_row_bitmap <= 16'b0000000000000000;
		15'h0a8d: char_row_bitmap <= 16'b0000000000000000;
		15'h0a8e: char_row_bitmap <= 16'b0111000000000000;
		15'h0a8f: char_row_bitmap <= 16'b0100100000000000;
		15'h0a90: char_row_bitmap <= 16'b0111000000000000;
		15'h0a91: char_row_bitmap <= 16'b0100100000000000;
		15'h0a92: char_row_bitmap <= 16'b0111000000000000;
		15'h0a93: char_row_bitmap <= 16'b0000000000000000;
		15'h0a94: char_row_bitmap <= 16'b0000001111000000;
		15'h0a95: char_row_bitmap <= 16'b0000001000000000;
		15'h0a96: char_row_bitmap <= 16'b0000001100000000;
		15'h0a97: char_row_bitmap <= 16'b0000001000000000;
		15'h0a98: char_row_bitmap <= 16'b0000001111000000;
		15'h0a99: char_row_bitmap <= 16'b0000000000000000;
		15'h0a9a: char_row_bitmap <= 16'b0000000000010000;
		15'h0a9b: char_row_bitmap <= 16'b0000000000010000;
		15'h0a9c: char_row_bitmap <= 16'b0000000000010000;
		15'h0a9d: char_row_bitmap <= 16'b0000000000010000;
		15'h0a9e: char_row_bitmap <= 16'b0000000000011110;
		15'h0a9f: char_row_bitmap <= 16'b0000000000000000;
		15'h0aa0: char_row_bitmap <= 16'b0000000000000000;
		15'h0aa1: char_row_bitmap <= 16'b0000000000000000;
		15'h0aa2: char_row_bitmap <= 16'b0000000000000000;
		15'h0aa3: char_row_bitmap <= 16'b0000000000000000;
		15'h0aa4: char_row_bitmap <= 16'b0000000000000000;
		15'h0aa5: char_row_bitmap <= 16'b0001110000000000;
		15'h0aa6: char_row_bitmap <= 16'b0001001000000000;
		15'h0aa7: char_row_bitmap <= 16'b0001110000000000;
		15'h0aa8: char_row_bitmap <= 16'b0001001000000000;
		15'h0aa9: char_row_bitmap <= 16'b0001110000000000;
		15'h0aaa: char_row_bitmap <= 16'b0000000000000000;
		15'h0aab: char_row_bitmap <= 16'b0000000001110000;
		15'h0aac: char_row_bitmap <= 16'b0000000010000000;
		15'h0aad: char_row_bitmap <= 16'b0000000001100000;
		15'h0aae: char_row_bitmap <= 16'b0000000000010000;
		15'h0aaf: char_row_bitmap <= 16'b0000000011100000;
		15'h0ab0: char_row_bitmap <= 16'b0000000000000000;
		15'h0ab1: char_row_bitmap <= 16'b0000000000000000;
		15'h0ab2: char_row_bitmap <= 16'b0000000000000000;
		15'h0ab3: char_row_bitmap <= 16'b0000000000000000;
		15'h0ab4: char_row_bitmap <= 16'b0000000000000000;
		15'h0ab5: char_row_bitmap <= 16'b0000000000000000;
		15'h0ab6: char_row_bitmap <= 16'b0111000000000000;
		15'h0ab7: char_row_bitmap <= 16'b0010000000000000;
		15'h0ab8: char_row_bitmap <= 16'b0010000000000000;
		15'h0ab9: char_row_bitmap <= 16'b0010000000000000;
		15'h0aba: char_row_bitmap <= 16'b0010000000000000;
		15'h0abb: char_row_bitmap <= 16'b0000000000000000;
		15'h0abc: char_row_bitmap <= 16'b0000001100000000;
		15'h0abd: char_row_bitmap <= 16'b0000010010000000;
		15'h0abe: char_row_bitmap <= 16'b0000011110000000;
		15'h0abf: char_row_bitmap <= 16'b0000010010000000;
		15'h0ac0: char_row_bitmap <= 16'b0000010010000000;
		15'h0ac1: char_row_bitmap <= 16'b0000000000000000;
		15'h0ac2: char_row_bitmap <= 16'b0000000000111000;
		15'h0ac3: char_row_bitmap <= 16'b0000000000100100;
		15'h0ac4: char_row_bitmap <= 16'b0000000000111000;
		15'h0ac5: char_row_bitmap <= 16'b0000000000100100;
		15'h0ac6: char_row_bitmap <= 16'b0000000000111000;
		15'h0ac7: char_row_bitmap <= 16'b0000000000000000;
		15'h0ac8: char_row_bitmap <= 16'b0000000000000000;
		15'h0ac9: char_row_bitmap <= 16'b0000000000000000;
		15'h0aca: char_row_bitmap <= 16'b0000000000000000;
		15'h0acb: char_row_bitmap <= 16'b0000000000000000;
		15'h0acc: char_row_bitmap <= 16'b0000000000000000;
		15'h0acd: char_row_bitmap <= 16'b0001000000000000;
		15'h0ace: char_row_bitmap <= 16'b0001000000000000;
		15'h0acf: char_row_bitmap <= 16'b0001000000000000;
		15'h0ad0: char_row_bitmap <= 16'b0001000000000000;
		15'h0ad1: char_row_bitmap <= 16'b0001111000000000;
		15'h0ad2: char_row_bitmap <= 16'b0000000000000000;
		15'h0ad3: char_row_bitmap <= 16'b0000000011110000;
		15'h0ad4: char_row_bitmap <= 16'b0000000010000000;
		15'h0ad5: char_row_bitmap <= 16'b0000000011000000;
		15'h0ad6: char_row_bitmap <= 16'b0000000010000000;
		15'h0ad7: char_row_bitmap <= 16'b0000000010000000;
		15'h0ad8: char_row_bitmap <= 16'b0000000000000000;
		15'h0ad9: char_row_bitmap <= 16'b0000000000000000;
		15'h0ada: char_row_bitmap <= 16'b0000000000000000;
		15'h0adb: char_row_bitmap <= 16'b0000000000000000;
		15'h0adc: char_row_bitmap <= 16'b0000000000000000;
		15'h0add: char_row_bitmap <= 16'b0000000000000000;
		15'h0ade: char_row_bitmap <= 16'b0000000000000000;
		15'h0adf: char_row_bitmap <= 16'b0000000000000000;
		15'h0ae0: char_row_bitmap <= 16'b0000000000000000;
		15'h0ae1: char_row_bitmap <= 16'b0001000100000000;
		15'h0ae2: char_row_bitmap <= 16'b0001000100000000;
		15'h0ae3: char_row_bitmap <= 16'b0001000100000000;
		15'h0ae4: char_row_bitmap <= 16'b0000101000000000;
		15'h0ae5: char_row_bitmap <= 16'b0000010000000000;
		15'h0ae6: char_row_bitmap <= 16'b0000000000000000;
		15'h0ae7: char_row_bitmap <= 16'b0000000001110000;
		15'h0ae8: char_row_bitmap <= 16'b0000000000100000;
		15'h0ae9: char_row_bitmap <= 16'b0000000000100000;
		15'h0aea: char_row_bitmap <= 16'b0000000000100000;
		15'h0aeb: char_row_bitmap <= 16'b0000000000100000;
		15'h0aec: char_row_bitmap <= 16'b0000000000000000;
		15'h0aed: char_row_bitmap <= 16'b0000000000000000;
		15'h0aee: char_row_bitmap <= 16'b0000000000000000;
		15'h0aef: char_row_bitmap <= 16'b0000000000000000;
		15'h0af0: char_row_bitmap <= 16'b0000000000000000;
		15'h0af1: char_row_bitmap <= 16'b0000000000000000;
		15'h0af2: char_row_bitmap <= 16'b0000000000000000;
		15'h0af3: char_row_bitmap <= 16'b0000000000000000;
		15'h0af4: char_row_bitmap <= 16'b0000000000000000;
		15'h0af5: char_row_bitmap <= 16'b0001111000000000;
		15'h0af6: char_row_bitmap <= 16'b0001000000000000;
		15'h0af7: char_row_bitmap <= 16'b0001100000000000;
		15'h0af8: char_row_bitmap <= 16'b0001000000000000;
		15'h0af9: char_row_bitmap <= 16'b0001000000000000;
		15'h0afa: char_row_bitmap <= 16'b0000000000000000;
		15'h0afb: char_row_bitmap <= 16'b0000000011110000;
		15'h0afc: char_row_bitmap <= 16'b0000000010000000;
		15'h0afd: char_row_bitmap <= 16'b0000000011000000;
		15'h0afe: char_row_bitmap <= 16'b0000000010000000;
		15'h0aff: char_row_bitmap <= 16'b0000000010000000;
		15'h0b00: char_row_bitmap <= 16'b0000000000000000;
		15'h0b01: char_row_bitmap <= 16'b0000000000000000;
		15'h0b02: char_row_bitmap <= 16'b0000000000000000;
		15'h0b03: char_row_bitmap <= 16'b0000000000000000;
		15'h0b04: char_row_bitmap <= 16'b0000000000000000;
		15'h0b05: char_row_bitmap <= 16'b0000000000000000;
		15'h0b06: char_row_bitmap <= 16'b0000000000000000;
		15'h0b07: char_row_bitmap <= 16'b0000000000000000;
		15'h0b08: char_row_bitmap <= 16'b0000000000000000;
		15'h0b09: char_row_bitmap <= 16'b0000111000000000;
		15'h0b0a: char_row_bitmap <= 16'b0001000000000000;
		15'h0b0b: char_row_bitmap <= 16'b0001000000000000;
		15'h0b0c: char_row_bitmap <= 16'b0001000000000000;
		15'h0b0d: char_row_bitmap <= 16'b0000111000000000;
		15'h0b0e: char_row_bitmap <= 16'b0000000000000000;
		15'h0b0f: char_row_bitmap <= 16'b0000000011100000;
		15'h0b10: char_row_bitmap <= 16'b0000000010010000;
		15'h0b11: char_row_bitmap <= 16'b0000000011100000;
		15'h0b12: char_row_bitmap <= 16'b0000000010100000;
		15'h0b13: char_row_bitmap <= 16'b0000000010010000;
		15'h0b14: char_row_bitmap <= 16'b0000000000000000;
		15'h0b15: char_row_bitmap <= 16'b0000000000000000;
		15'h0b16: char_row_bitmap <= 16'b0000000000000000;
		15'h0b17: char_row_bitmap <= 16'b0000000000000000;
		15'h0b18: char_row_bitmap <= 16'b0000000000000000;
		15'h0b19: char_row_bitmap <= 16'b0000000000000000;
		15'h0b1a: char_row_bitmap <= 16'b0000000000000000;
		15'h0b1b: char_row_bitmap <= 16'b0000000000000000;
		15'h0b1c: char_row_bitmap <= 16'b0000000000000000;
		15'h0b1d: char_row_bitmap <= 16'b0000111000000000;
		15'h0b1e: char_row_bitmap <= 16'b0001000000000000;
		15'h0b1f: char_row_bitmap <= 16'b0000110000000000;
		15'h0b20: char_row_bitmap <= 16'b0000001000000000;
		15'h0b21: char_row_bitmap <= 16'b0001110000000000;
		15'h0b22: char_row_bitmap <= 16'b0000000000000000;
		15'h0b23: char_row_bitmap <= 16'b0000000001110000;
		15'h0b24: char_row_bitmap <= 16'b0000000010000000;
		15'h0b25: char_row_bitmap <= 16'b0000000001100000;
		15'h0b26: char_row_bitmap <= 16'b0000000000010000;
		15'h0b27: char_row_bitmap <= 16'b0000000011100000;
		15'h0b28: char_row_bitmap <= 16'b0000000000000000;
		15'h0b29: char_row_bitmap <= 16'b0000000000000000;
		15'h0b2a: char_row_bitmap <= 16'b0000000000000000;
		15'h0b2b: char_row_bitmap <= 16'b0000000000000000;
		15'h0b2c: char_row_bitmap <= 16'b0000000000000000;
		15'h0b2d: char_row_bitmap <= 16'b0000000000000000;
		15'h0b2e: char_row_bitmap <= 16'b0000000000000000;
		15'h0b2f: char_row_bitmap <= 16'b0000000000000000;
		15'h0b30: char_row_bitmap <= 16'b0000000000000000;
		15'h0b31: char_row_bitmap <= 16'b0000111000000000;
		15'h0b32: char_row_bitmap <= 16'b0001000000000000;
		15'h0b33: char_row_bitmap <= 16'b0000110000000000;
		15'h0b34: char_row_bitmap <= 16'b0000001000000000;
		15'h0b35: char_row_bitmap <= 16'b0001110000000000;
		15'h0b36: char_row_bitmap <= 16'b0000000000000000;
		15'h0b37: char_row_bitmap <= 16'b0000000011100000;
		15'h0b38: char_row_bitmap <= 16'b0000000001000000;
		15'h0b39: char_row_bitmap <= 16'b0000000001000000;
		15'h0b3a: char_row_bitmap <= 16'b0000000001000000;
		15'h0b3b: char_row_bitmap <= 16'b0000000011100000;
		15'h0b3c: char_row_bitmap <= 16'b0000000000000000;
		15'h0b3d: char_row_bitmap <= 16'b0000000000000000;
		15'h0b3e: char_row_bitmap <= 16'b0000000000000000;
		15'h0b3f: char_row_bitmap <= 16'b0000000000000000;
		15'h0b40: char_row_bitmap <= 16'b0000000000000000;
		15'h0b41: char_row_bitmap <= 16'b0000000000000000;
		15'h0b42: char_row_bitmap <= 16'b0111000000000000;
		15'h0b43: char_row_bitmap <= 16'b0100100000000000;
		15'h0b44: char_row_bitmap <= 16'b0100100000000000;
		15'h0b45: char_row_bitmap <= 16'b0100100000000000;
		15'h0b46: char_row_bitmap <= 16'b0111000000000000;
		15'h0b47: char_row_bitmap <= 16'b0000000000000000;
		15'h0b48: char_row_bitmap <= 16'b0000001000000000;
		15'h0b49: char_row_bitmap <= 16'b0000001000000000;
		15'h0b4a: char_row_bitmap <= 16'b0000001000000000;
		15'h0b4b: char_row_bitmap <= 16'b0000001000000000;
		15'h0b4c: char_row_bitmap <= 16'b0000001111000000;
		15'h0b4d: char_row_bitmap <= 16'b0000000000000000;
		15'h0b4e: char_row_bitmap <= 16'b0000000000011110;
		15'h0b4f: char_row_bitmap <= 16'b0000000000010000;
		15'h0b50: char_row_bitmap <= 16'b0000000000011000;
		15'h0b51: char_row_bitmap <= 16'b0000000000010000;
		15'h0b52: char_row_bitmap <= 16'b0000000000011110;
		15'h0b53: char_row_bitmap <= 16'b0000000000000000;
		15'h0b54: char_row_bitmap <= 16'b0000000000000000;
		15'h0b55: char_row_bitmap <= 16'b0000000000000000;
		15'h0b56: char_row_bitmap <= 16'b0111000000000000;
		15'h0b57: char_row_bitmap <= 16'b0100100000000000;
		15'h0b58: char_row_bitmap <= 16'b0100100000000000;
		15'h0b59: char_row_bitmap <= 16'b0100100000000000;
		15'h0b5a: char_row_bitmap <= 16'b0111000000000000;
		15'h0b5b: char_row_bitmap <= 16'b0000000000000000;
		15'h0b5c: char_row_bitmap <= 16'b0000000111000000;
		15'h0b5d: char_row_bitmap <= 16'b0000001000000000;
		15'h0b5e: char_row_bitmap <= 16'b0000001000000000;
		15'h0b5f: char_row_bitmap <= 16'b0000001000000000;
		15'h0b60: char_row_bitmap <= 16'b0000000111000000;
		15'h0b61: char_row_bitmap <= 16'b0000000000000000;
		15'h0b62: char_row_bitmap <= 16'b0000000000001000;
		15'h0b63: char_row_bitmap <= 16'b0000000000011000;
		15'h0b64: char_row_bitmap <= 16'b0000000000001000;
		15'h0b65: char_row_bitmap <= 16'b0000000000001000;
		15'h0b66: char_row_bitmap <= 16'b0000000000011100;
		15'h0b67: char_row_bitmap <= 16'b0000000000000000;
		15'h0b68: char_row_bitmap <= 16'b0000000000000000;
		15'h0b69: char_row_bitmap <= 16'b0000000000000000;
		15'h0b6a: char_row_bitmap <= 16'b0111000000000000;
		15'h0b6b: char_row_bitmap <= 16'b0100100000000000;
		15'h0b6c: char_row_bitmap <= 16'b0100100000000000;
		15'h0b6d: char_row_bitmap <= 16'b0100100000000000;
		15'h0b6e: char_row_bitmap <= 16'b0111000000000000;
		15'h0b6f: char_row_bitmap <= 16'b0000000000000000;
		15'h0b70: char_row_bitmap <= 16'b0000000111000000;
		15'h0b71: char_row_bitmap <= 16'b0000001000000000;
		15'h0b72: char_row_bitmap <= 16'b0000001000000000;
		15'h0b73: char_row_bitmap <= 16'b0000001000000000;
		15'h0b74: char_row_bitmap <= 16'b0000000111000000;
		15'h0b75: char_row_bitmap <= 16'b0000000000000000;
		15'h0b76: char_row_bitmap <= 16'b0000000000011000;
		15'h0b77: char_row_bitmap <= 16'b0000000000000100;
		15'h0b78: char_row_bitmap <= 16'b0000000000001000;
		15'h0b79: char_row_bitmap <= 16'b0000000000010000;
		15'h0b7a: char_row_bitmap <= 16'b0000000000011100;
		15'h0b7b: char_row_bitmap <= 16'b0000000000000000;
		15'h0b7c: char_row_bitmap <= 16'b0000000000000000;
		15'h0b7d: char_row_bitmap <= 16'b0000000000000000;
		15'h0b7e: char_row_bitmap <= 16'b0111000000000000;
		15'h0b7f: char_row_bitmap <= 16'b0100100000000000;
		15'h0b80: char_row_bitmap <= 16'b0100100000000000;
		15'h0b81: char_row_bitmap <= 16'b0100100000000000;
		15'h0b82: char_row_bitmap <= 16'b0111000000000000;
		15'h0b83: char_row_bitmap <= 16'b0000000000000000;
		15'h0b84: char_row_bitmap <= 16'b0000000111000000;
		15'h0b85: char_row_bitmap <= 16'b0000001000000000;
		15'h0b86: char_row_bitmap <= 16'b0000001000000000;
		15'h0b87: char_row_bitmap <= 16'b0000001000000000;
		15'h0b88: char_row_bitmap <= 16'b0000000111000000;
		15'h0b89: char_row_bitmap <= 16'b0000000000000000;
		15'h0b8a: char_row_bitmap <= 16'b0000000000011000;
		15'h0b8b: char_row_bitmap <= 16'b0000000000000100;
		15'h0b8c: char_row_bitmap <= 16'b0000000000001000;
		15'h0b8d: char_row_bitmap <= 16'b0000000000000100;
		15'h0b8e: char_row_bitmap <= 16'b0000000000011000;
		15'h0b8f: char_row_bitmap <= 16'b0000000000000000;
		15'h0b90: char_row_bitmap <= 16'b0000000000000000;
		15'h0b91: char_row_bitmap <= 16'b0000000000000000;
		15'h0b92: char_row_bitmap <= 16'b0111000000000000;
		15'h0b93: char_row_bitmap <= 16'b0100100000000000;
		15'h0b94: char_row_bitmap <= 16'b0100100000000000;
		15'h0b95: char_row_bitmap <= 16'b0100100000000000;
		15'h0b96: char_row_bitmap <= 16'b0111000000000000;
		15'h0b97: char_row_bitmap <= 16'b0000000000000000;
		15'h0b98: char_row_bitmap <= 16'b0000000111000000;
		15'h0b99: char_row_bitmap <= 16'b0000001000000000;
		15'h0b9a: char_row_bitmap <= 16'b0000001000000000;
		15'h0b9b: char_row_bitmap <= 16'b0000001000000000;
		15'h0b9c: char_row_bitmap <= 16'b0000000111000000;
		15'h0b9d: char_row_bitmap <= 16'b0000000000000000;
		15'h0b9e: char_row_bitmap <= 16'b0000000000010100;
		15'h0b9f: char_row_bitmap <= 16'b0000000000010100;
		15'h0ba0: char_row_bitmap <= 16'b0000000000011100;
		15'h0ba1: char_row_bitmap <= 16'b0000000000000100;
		15'h0ba2: char_row_bitmap <= 16'b0000000000000100;
		15'h0ba3: char_row_bitmap <= 16'b0000000000000000;
		15'h0ba4: char_row_bitmap <= 16'b0000000000000000;
		15'h0ba5: char_row_bitmap <= 16'b0000000000000000;
		15'h0ba6: char_row_bitmap <= 16'b0100100000000000;
		15'h0ba7: char_row_bitmap <= 16'b0110100000000000;
		15'h0ba8: char_row_bitmap <= 16'b0101100000000000;
		15'h0ba9: char_row_bitmap <= 16'b0100100000000000;
		15'h0baa: char_row_bitmap <= 16'b0100100000000000;
		15'h0bab: char_row_bitmap <= 16'b0000000000000000;
		15'h0bac: char_row_bitmap <= 16'b0000000110000000;
		15'h0bad: char_row_bitmap <= 16'b0000001001000000;
		15'h0bae: char_row_bitmap <= 16'b0000001111000000;
		15'h0baf: char_row_bitmap <= 16'b0000001001000000;
		15'h0bb0: char_row_bitmap <= 16'b0000001001000000;
		15'h0bb1: char_row_bitmap <= 16'b0000000000000000;
		15'h0bb2: char_row_bitmap <= 16'b0000000000010010;
		15'h0bb3: char_row_bitmap <= 16'b0000000000010100;
		15'h0bb4: char_row_bitmap <= 16'b0000000000011000;
		15'h0bb5: char_row_bitmap <= 16'b0000000000010100;
		15'h0bb6: char_row_bitmap <= 16'b0000000000010010;
		15'h0bb7: char_row_bitmap <= 16'b0000000000000000;
		15'h0bb8: char_row_bitmap <= 16'b0000000000000000;
		15'h0bb9: char_row_bitmap <= 16'b0000000000000000;
		15'h0bba: char_row_bitmap <= 16'b0011100000000000;
		15'h0bbb: char_row_bitmap <= 16'b0100000000000000;
		15'h0bbc: char_row_bitmap <= 16'b0011000000000000;
		15'h0bbd: char_row_bitmap <= 16'b0000100000000000;
		15'h0bbe: char_row_bitmap <= 16'b0111000000000000;
		15'h0bbf: char_row_bitmap <= 16'b0000000000000000;
		15'h0bc0: char_row_bitmap <= 16'b0000001010000000;
		15'h0bc1: char_row_bitmap <= 16'b0000001010000000;
		15'h0bc2: char_row_bitmap <= 16'b0000000100000000;
		15'h0bc3: char_row_bitmap <= 16'b0000000100000000;
		15'h0bc4: char_row_bitmap <= 16'b0000000100000000;
		15'h0bc5: char_row_bitmap <= 16'b0000000000000000;
		15'h0bc6: char_row_bitmap <= 16'b0000000000100100;
		15'h0bc7: char_row_bitmap <= 16'b0000000000110100;
		15'h0bc8: char_row_bitmap <= 16'b0000000000101100;
		15'h0bc9: char_row_bitmap <= 16'b0000000000100100;
		15'h0bca: char_row_bitmap <= 16'b0000000000100100;
		15'h0bcb: char_row_bitmap <= 16'b0000000000000000;
		15'h0bcc: char_row_bitmap <= 16'b0000000000000000;
		15'h0bcd: char_row_bitmap <= 16'b0000000000000000;
		15'h0bce: char_row_bitmap <= 16'b0111100000000000;
		15'h0bcf: char_row_bitmap <= 16'b0100000000000000;
		15'h0bd0: char_row_bitmap <= 16'b0110000000000000;
		15'h0bd1: char_row_bitmap <= 16'b0100000000000000;
		15'h0bd2: char_row_bitmap <= 16'b0111100000000000;
		15'h0bd3: char_row_bitmap <= 16'b0000000000000000;
		15'h0bd4: char_row_bitmap <= 16'b0000001110000000;
		15'h0bd5: char_row_bitmap <= 16'b0000000100000000;
		15'h0bd6: char_row_bitmap <= 16'b0000000100000000;
		15'h0bd7: char_row_bitmap <= 16'b0000000100000000;
		15'h0bd8: char_row_bitmap <= 16'b0000000100000000;
		15'h0bd9: char_row_bitmap <= 16'b0000000000000000;
		15'h0bda: char_row_bitmap <= 16'b0000000000011100;
		15'h0bdb: char_row_bitmap <= 16'b0000000000010010;
		15'h0bdc: char_row_bitmap <= 16'b0000000000011100;
		15'h0bdd: char_row_bitmap <= 16'b0000000000010010;
		15'h0bde: char_row_bitmap <= 16'b0000000000011100;
		15'h0bdf: char_row_bitmap <= 16'b0000000000000000;
		15'h0be0: char_row_bitmap <= 16'b0000000000000000;
		15'h0be1: char_row_bitmap <= 16'b0000000000000000;
		15'h0be2: char_row_bitmap <= 16'b0011100000000000;
		15'h0be3: char_row_bitmap <= 16'b0100000000000000;
		15'h0be4: char_row_bitmap <= 16'b0100000000000000;
		15'h0be5: char_row_bitmap <= 16'b0100000000000000;
		15'h0be6: char_row_bitmap <= 16'b0011100000000000;
		15'h0be7: char_row_bitmap <= 16'b0000000000000000;
		15'h0be8: char_row_bitmap <= 16'b0000000110000000;
		15'h0be9: char_row_bitmap <= 16'b0000001001000000;
		15'h0bea: char_row_bitmap <= 16'b0000001111000000;
		15'h0beb: char_row_bitmap <= 16'b0000001001000000;
		15'h0bec: char_row_bitmap <= 16'b0000001001000000;
		15'h0bed: char_row_bitmap <= 16'b0000000000000000;
		15'h0bee: char_row_bitmap <= 16'b0000000000010010;
		15'h0bef: char_row_bitmap <= 16'b0000000000011010;
		15'h0bf0: char_row_bitmap <= 16'b0000000000010110;
		15'h0bf1: char_row_bitmap <= 16'b0000000000010010;
		15'h0bf2: char_row_bitmap <= 16'b0000000000010010;
		15'h0bf3: char_row_bitmap <= 16'b0000000000000000;
		15'h0bf4: char_row_bitmap <= 16'b0000000000000000;
		15'h0bf5: char_row_bitmap <= 16'b0000000000000000;
		15'h0bf6: char_row_bitmap <= 16'b0000000000000000;
		15'h0bf7: char_row_bitmap <= 16'b0000000000000000;
		15'h0bf8: char_row_bitmap <= 16'b0000000000000000;
		15'h0bf9: char_row_bitmap <= 16'b0001111000000000;
		15'h0bfa: char_row_bitmap <= 16'b0001000000000000;
		15'h0bfb: char_row_bitmap <= 16'b0001100000000000;
		15'h0bfc: char_row_bitmap <= 16'b0001000000000000;
		15'h0bfd: char_row_bitmap <= 16'b0001111000000000;
		15'h0bfe: char_row_bitmap <= 16'b0000000000000000;
		15'h0bff: char_row_bitmap <= 16'b0000000010001000;
		15'h0c00: char_row_bitmap <= 16'b0000000011011000;
		15'h0c01: char_row_bitmap <= 16'b0000000010101000;
		15'h0c02: char_row_bitmap <= 16'b0000000010001000;
		15'h0c03: char_row_bitmap <= 16'b0000000010001000;
		15'h0c04: char_row_bitmap <= 16'b0000000000000000;
		15'h0c05: char_row_bitmap <= 16'b0000000000000000;
		15'h0c06: char_row_bitmap <= 16'b0000000000000000;
		15'h0c07: char_row_bitmap <= 16'b0000000000000000;
		15'h0c08: char_row_bitmap <= 16'b0000000000000000;
		15'h0c09: char_row_bitmap <= 16'b0000000000000000;
		15'h0c0a: char_row_bitmap <= 16'b0011100000000000;
		15'h0c0b: char_row_bitmap <= 16'b0100000000000000;
		15'h0c0c: char_row_bitmap <= 16'b0011000000000000;
		15'h0c0d: char_row_bitmap <= 16'b0000100000000000;
		15'h0c0e: char_row_bitmap <= 16'b0111000000000000;
		15'h0c0f: char_row_bitmap <= 16'b0000000000000000;
		15'h0c10: char_row_bitmap <= 16'b0000001001000000;
		15'h0c11: char_row_bitmap <= 16'b0000001001000000;
		15'h0c12: char_row_bitmap <= 16'b0000001001000000;
		15'h0c13: char_row_bitmap <= 16'b0000001001000000;
		15'h0c14: char_row_bitmap <= 16'b0000000110000000;
		15'h0c15: char_row_bitmap <= 16'b0000000000000000;
		15'h0c16: char_row_bitmap <= 16'b0000000000011100;
		15'h0c17: char_row_bitmap <= 16'b0000000000010010;
		15'h0c18: char_row_bitmap <= 16'b0000000000011100;
		15'h0c19: char_row_bitmap <= 16'b0000000000010010;
		15'h0c1a: char_row_bitmap <= 16'b0000000000011100;
		15'h0c1b: char_row_bitmap <= 16'b0000000000000000;
		15'h0c1c: char_row_bitmap <= 16'b0000000000000000;
		15'h0c1d: char_row_bitmap <= 16'b0000000000000000;
		15'h0c1e: char_row_bitmap <= 16'b0111100000000000;
		15'h0c1f: char_row_bitmap <= 16'b0100000000000000;
		15'h0c20: char_row_bitmap <= 16'b0110000000000000;
		15'h0c21: char_row_bitmap <= 16'b0100000000000000;
		15'h0c22: char_row_bitmap <= 16'b0111100000000000;
		15'h0c23: char_row_bitmap <= 16'b0000000000000000;
		15'h0c24: char_row_bitmap <= 16'b0000000111000000;
		15'h0c25: char_row_bitmap <= 16'b0000001000000000;
		15'h0c26: char_row_bitmap <= 16'b0000000110000000;
		15'h0c27: char_row_bitmap <= 16'b0000000001000000;
		15'h0c28: char_row_bitmap <= 16'b0000001110000000;
		15'h0c29: char_row_bitmap <= 16'b0000000000000000;
		15'h0c2a: char_row_bitmap <= 16'b0000000000001110;
		15'h0c2b: char_row_bitmap <= 16'b0000000000010000;
		15'h0c2c: char_row_bitmap <= 16'b0000000000010000;
		15'h0c2d: char_row_bitmap <= 16'b0000000000010000;
		15'h0c2e: char_row_bitmap <= 16'b0000000000001110;
		15'h0c2f: char_row_bitmap <= 16'b0000000000000000;
		15'h0c30: char_row_bitmap <= 16'b0000000000000000;
		15'h0c31: char_row_bitmap <= 16'b0000000000000000;
		15'h0c32: char_row_bitmap <= 16'b0000000000000000;
		15'h0c33: char_row_bitmap <= 16'b0000000000000000;
		15'h0c34: char_row_bitmap <= 16'b0000000000000000;
		15'h0c35: char_row_bitmap <= 16'b0001111000000000;
		15'h0c36: char_row_bitmap <= 16'b0001000000000000;
		15'h0c37: char_row_bitmap <= 16'b0001100000000000;
		15'h0c38: char_row_bitmap <= 16'b0001000000000000;
		15'h0c39: char_row_bitmap <= 16'b0001000000000000;
		15'h0c3a: char_row_bitmap <= 16'b0000000000000000;
		15'h0c3b: char_row_bitmap <= 16'b0000000001110000;
		15'h0c3c: char_row_bitmap <= 16'b0000000010000000;
		15'h0c3d: char_row_bitmap <= 16'b0000000001100000;
		15'h0c3e: char_row_bitmap <= 16'b0000000000010000;
		15'h0c3f: char_row_bitmap <= 16'b0000000011100000;
		15'h0c40: char_row_bitmap <= 16'b0000000000000000;
		15'h0c41: char_row_bitmap <= 16'b0000000000000000;
		15'h0c42: char_row_bitmap <= 16'b0000000000000000;
		15'h0c43: char_row_bitmap <= 16'b0000000000000000;
		15'h0c44: char_row_bitmap <= 16'b0000000000000000;
		15'h0c45: char_row_bitmap <= 16'b0000000000000000;
		15'h0c46: char_row_bitmap <= 16'b0000000000000000;
		15'h0c47: char_row_bitmap <= 16'b0000000000000000;
		15'h0c48: char_row_bitmap <= 16'b0000000000000000;
		15'h0c49: char_row_bitmap <= 16'b0000110000000000;
		15'h0c4a: char_row_bitmap <= 16'b0001000000000000;
		15'h0c4b: char_row_bitmap <= 16'b0001011000000000;
		15'h0c4c: char_row_bitmap <= 16'b0001001000000000;
		15'h0c4d: char_row_bitmap <= 16'b0000111000000000;
		15'h0c4e: char_row_bitmap <= 16'b0000000000000000;
		15'h0c4f: char_row_bitmap <= 16'b0000000001110000;
		15'h0c50: char_row_bitmap <= 16'b0000000010000000;
		15'h0c51: char_row_bitmap <= 16'b0000000001100000;
		15'h0c52: char_row_bitmap <= 16'b0000000000010000;
		15'h0c53: char_row_bitmap <= 16'b0000000011100000;
		15'h0c54: char_row_bitmap <= 16'b0000000000000000;
		15'h0c55: char_row_bitmap <= 16'b0000000000000000;
		15'h0c56: char_row_bitmap <= 16'b0000000000000000;
		15'h0c57: char_row_bitmap <= 16'b0000000000000000;
		15'h0c58: char_row_bitmap <= 16'b0000000000000000;
		15'h0c59: char_row_bitmap <= 16'b0000000000000000;
		15'h0c5a: char_row_bitmap <= 16'b0000000000000000;
		15'h0c5b: char_row_bitmap <= 16'b0000000000000000;
		15'h0c5c: char_row_bitmap <= 16'b0000000000000000;
		15'h0c5d: char_row_bitmap <= 16'b0001110000000000;
		15'h0c5e: char_row_bitmap <= 16'b0001001000000000;
		15'h0c5f: char_row_bitmap <= 16'b0001110000000000;
		15'h0c60: char_row_bitmap <= 16'b0001010000000000;
		15'h0c61: char_row_bitmap <= 16'b0001001000000000;
		15'h0c62: char_row_bitmap <= 16'b0000000000000000;
		15'h0c63: char_row_bitmap <= 16'b0000000001110000;
		15'h0c64: char_row_bitmap <= 16'b0000000010000000;
		15'h0c65: char_row_bitmap <= 16'b0000000001100000;
		15'h0c66: char_row_bitmap <= 16'b0000000000010000;
		15'h0c67: char_row_bitmap <= 16'b0000000011100000;
		15'h0c68: char_row_bitmap <= 16'b0000000000000000;
		15'h0c69: char_row_bitmap <= 16'b0000000000000000;
		15'h0c6a: char_row_bitmap <= 16'b0000000000000000;
		15'h0c6b: char_row_bitmap <= 16'b0000000000000000;
		15'h0c6c: char_row_bitmap <= 16'b0000000000000000;
		15'h0c6d: char_row_bitmap <= 16'b0000000000000000;
		15'h0c6e: char_row_bitmap <= 16'b0000000000000000;
		15'h0c6f: char_row_bitmap <= 16'b0000000000000000;
		15'h0c70: char_row_bitmap <= 16'b0000000000000000;
		15'h0c71: char_row_bitmap <= 16'b0001001000000000;
		15'h0c72: char_row_bitmap <= 16'b0001001000000000;
		15'h0c73: char_row_bitmap <= 16'b0001001000000000;
		15'h0c74: char_row_bitmap <= 16'b0001001000000000;
		15'h0c75: char_row_bitmap <= 16'b0000110000000000;
		15'h0c76: char_row_bitmap <= 16'b0000000000000000;
		15'h0c77: char_row_bitmap <= 16'b0000000001110000;
		15'h0c78: char_row_bitmap <= 16'b0000000010000000;
		15'h0c79: char_row_bitmap <= 16'b0000000001100000;
		15'h0c7a: char_row_bitmap <= 16'b0000000000010000;
		15'h0c7b: char_row_bitmap <= 16'b0000000011100000;
		15'h0c7c: char_row_bitmap <= 16'b0000000000000000;
		15'h0c7d: char_row_bitmap <= 16'b0000000000000000;
		15'h0c7e: char_row_bitmap <= 16'b0000000000000000;
		15'h0c7f: char_row_bitmap <= 16'b0000000000000000;
		15'h0c80: char_row_bitmap <= 16'b0000000000000000;
		15'h0c81: char_row_bitmap <= 16'b0000000000000000;
		15'h0c82: char_row_bitmap <= 16'b0000000000000000;
		15'h0c83: char_row_bitmap <= 16'b0000000000000000;
		15'h0c84: char_row_bitmap <= 16'b0000000000000000;
		15'h0c85: char_row_bitmap <= 16'b0000000000000000;
		15'h0c86: char_row_bitmap <= 16'b0000111000011000;
		15'h0c87: char_row_bitmap <= 16'b0001111100110000;
		15'h0c88: char_row_bitmap <= 16'b0011101110110000;
		15'h0c89: char_row_bitmap <= 16'b0011000111100000;
		15'h0c8a: char_row_bitmap <= 16'b0011000011100000;
		15'h0c8b: char_row_bitmap <= 16'b0011000011100000;
		15'h0c8c: char_row_bitmap <= 16'b0011000111100000;
		15'h0c8d: char_row_bitmap <= 16'b0011101110110000;
		15'h0c8e: char_row_bitmap <= 16'b0001111100110000;
		15'h0c8f: char_row_bitmap <= 16'b0000111000011000;
		15'h0c90: char_row_bitmap <= 16'b0000000000000000;
		15'h0c91: char_row_bitmap <= 16'b0000000000000000;
		15'h0c92: char_row_bitmap <= 16'b0000000000000000;
		15'h0c93: char_row_bitmap <= 16'b0000000000000000;
		15'h0c94: char_row_bitmap <= 16'b0000000000000000;
		15'h0c95: char_row_bitmap <= 16'b0000000000000000;
		15'h0c96: char_row_bitmap <= 16'b0000001100000000;
		15'h0c97: char_row_bitmap <= 16'b0000011110000000;
		15'h0c98: char_row_bitmap <= 16'b0000111011000000;
		15'h0c99: char_row_bitmap <= 16'b0000110011000000;
		15'h0c9a: char_row_bitmap <= 16'b0001110111000000;
		15'h0c9b: char_row_bitmap <= 16'b0001100110000000;
		15'h0c9c: char_row_bitmap <= 16'b0001111110000000;
		15'h0c9d: char_row_bitmap <= 16'b0001111111000000;
		15'h0c9e: char_row_bitmap <= 16'b0001100011100000;
		15'h0c9f: char_row_bitmap <= 16'b0001100001100000;
		15'h0ca0: char_row_bitmap <= 16'b0001100001100000;
		15'h0ca1: char_row_bitmap <= 16'b0001100011100000;
		15'h0ca2: char_row_bitmap <= 16'b0001111111000000;
		15'h0ca3: char_row_bitmap <= 16'b0001111110000000;
		15'h0ca4: char_row_bitmap <= 16'b0001100000000000;
		15'h0ca5: char_row_bitmap <= 16'b0001100000000000;
		15'h0ca6: char_row_bitmap <= 16'b0001100000000000;
		15'h0ca7: char_row_bitmap <= 16'b0000000000000000;
		15'h0ca8: char_row_bitmap <= 16'b0000000000000000;
		15'h0ca9: char_row_bitmap <= 16'b0000000000000000;
		15'h0caa: char_row_bitmap <= 16'b0000000000000000;
		15'h0cab: char_row_bitmap <= 16'b0011111111100000;
		15'h0cac: char_row_bitmap <= 16'b0011111111100000;
		15'h0cad: char_row_bitmap <= 16'b0011000001100000;
		15'h0cae: char_row_bitmap <= 16'b0011000001100000;
		15'h0caf: char_row_bitmap <= 16'b0011000000000000;
		15'h0cb0: char_row_bitmap <= 16'b0011000000000000;
		15'h0cb1: char_row_bitmap <= 16'b0011000000000000;
		15'h0cb2: char_row_bitmap <= 16'b0011000000000000;
		15'h0cb3: char_row_bitmap <= 16'b0011000000000000;
		15'h0cb4: char_row_bitmap <= 16'b0011000000000000;
		15'h0cb5: char_row_bitmap <= 16'b0011000000000000;
		15'h0cb6: char_row_bitmap <= 16'b0011000000000000;
		15'h0cb7: char_row_bitmap <= 16'b0011000000000000;
		15'h0cb8: char_row_bitmap <= 16'b0000000000000000;
		15'h0cb9: char_row_bitmap <= 16'b0000000000000000;
		15'h0cba: char_row_bitmap <= 16'b0000000000000000;
		15'h0cbb: char_row_bitmap <= 16'b0000000000000000;
		15'h0cbc: char_row_bitmap <= 16'b0000000000000000;
		15'h0cbd: char_row_bitmap <= 16'b0000000000000000;
		15'h0cbe: char_row_bitmap <= 16'b0000000000000000;
		15'h0cbf: char_row_bitmap <= 16'b0000000000000000;
		15'h0cc0: char_row_bitmap <= 16'b0000000000000000;
		15'h0cc1: char_row_bitmap <= 16'b0000000000000000;
		15'h0cc2: char_row_bitmap <= 16'b0000000000000000;
		15'h0cc3: char_row_bitmap <= 16'b0000000000000000;
		15'h0cc4: char_row_bitmap <= 16'b0011111111110000;
		15'h0cc5: char_row_bitmap <= 16'b0011111111110000;
		15'h0cc6: char_row_bitmap <= 16'b0000110011000000;
		15'h0cc7: char_row_bitmap <= 16'b0000110011000000;
		15'h0cc8: char_row_bitmap <= 16'b0000110011000000;
		15'h0cc9: char_row_bitmap <= 16'b0000110011100000;
		15'h0cca: char_row_bitmap <= 16'b0000110001110000;
		15'h0ccb: char_row_bitmap <= 16'b0000110000110000;
		15'h0ccc: char_row_bitmap <= 16'b0000000000000000;
		15'h0ccd: char_row_bitmap <= 16'b0000000000000000;
		15'h0cce: char_row_bitmap <= 16'b0000000000000000;
		15'h0ccf: char_row_bitmap <= 16'b0000000000000000;
		15'h0cd0: char_row_bitmap <= 16'b0000000000000000;
		15'h0cd1: char_row_bitmap <= 16'b0000000000000000;
		15'h0cd2: char_row_bitmap <= 16'b0011111111110000;
		15'h0cd3: char_row_bitmap <= 16'b0011111111110000;
		15'h0cd4: char_row_bitmap <= 16'b0011100000110000;
		15'h0cd5: char_row_bitmap <= 16'b0001110000110000;
		15'h0cd6: char_row_bitmap <= 16'b0000111000000000;
		15'h0cd7: char_row_bitmap <= 16'b0000011100000000;
		15'h0cd8: char_row_bitmap <= 16'b0000001110000000;
		15'h0cd9: char_row_bitmap <= 16'b0000001110000000;
		15'h0cda: char_row_bitmap <= 16'b0000011100000000;
		15'h0cdb: char_row_bitmap <= 16'b0000111000000000;
		15'h0cdc: char_row_bitmap <= 16'b0001110000110000;
		15'h0cdd: char_row_bitmap <= 16'b0011100000110000;
		15'h0cde: char_row_bitmap <= 16'b0011111111110000;
		15'h0cdf: char_row_bitmap <= 16'b0011111111110000;
		15'h0ce0: char_row_bitmap <= 16'b0000000000000000;
		15'h0ce1: char_row_bitmap <= 16'b0000000000000000;
		15'h0ce2: char_row_bitmap <= 16'b0000000000000000;
		15'h0ce3: char_row_bitmap <= 16'b0000000000000000;
		15'h0ce4: char_row_bitmap <= 16'b0000000000000000;
		15'h0ce5: char_row_bitmap <= 16'b0000000000000000;
		15'h0ce6: char_row_bitmap <= 16'b0000000000000000;
		15'h0ce7: char_row_bitmap <= 16'b0000000000000000;
		15'h0ce8: char_row_bitmap <= 16'b0000000000000000;
		15'h0ce9: char_row_bitmap <= 16'b0000000000000000;
		15'h0cea: char_row_bitmap <= 16'b0000111000011000;
		15'h0ceb: char_row_bitmap <= 16'b0001111100110000;
		15'h0cec: char_row_bitmap <= 16'b0011101111110000;
		15'h0ced: char_row_bitmap <= 16'b0011000111100000;
		15'h0cee: char_row_bitmap <= 16'b0011000110000000;
		15'h0cef: char_row_bitmap <= 16'b0011000110000000;
		15'h0cf0: char_row_bitmap <= 16'b0011001110000000;
		15'h0cf1: char_row_bitmap <= 16'b0011101100000000;
		15'h0cf2: char_row_bitmap <= 16'b0001111100000000;
		15'h0cf3: char_row_bitmap <= 16'b0000111000000000;
		15'h0cf4: char_row_bitmap <= 16'b0000000000000000;
		15'h0cf5: char_row_bitmap <= 16'b0000000000000000;
		15'h0cf6: char_row_bitmap <= 16'b0000000000000000;
		15'h0cf7: char_row_bitmap <= 16'b0000000000000000;
		15'h0cf8: char_row_bitmap <= 16'b0000000000000000;
		15'h0cf9: char_row_bitmap <= 16'b0000000000000000;
		15'h0cfa: char_row_bitmap <= 16'b0000000000000000;
		15'h0cfb: char_row_bitmap <= 16'b0000000000000000;
		15'h0cfc: char_row_bitmap <= 16'b0000000000000000;
		15'h0cfd: char_row_bitmap <= 16'b0000000000000000;
		15'h0cfe: char_row_bitmap <= 16'b0001100001100000;
		15'h0cff: char_row_bitmap <= 16'b0001100001100000;
		15'h0d00: char_row_bitmap <= 16'b0001100001100000;
		15'h0d01: char_row_bitmap <= 16'b0001100001100000;
		15'h0d02: char_row_bitmap <= 16'b0001100001100000;
		15'h0d03: char_row_bitmap <= 16'b0001110011100000;
		15'h0d04: char_row_bitmap <= 16'b0001111111000000;
		15'h0d05: char_row_bitmap <= 16'b0001101110000000;
		15'h0d06: char_row_bitmap <= 16'b0001100000000000;
		15'h0d07: char_row_bitmap <= 16'b0001100000000000;
		15'h0d08: char_row_bitmap <= 16'b0011000000000000;
		15'h0d09: char_row_bitmap <= 16'b0011000000000000;
		15'h0d0a: char_row_bitmap <= 16'b0011000000000000;
		15'h0d0b: char_row_bitmap <= 16'b0011000000000000;
		15'h0d0c: char_row_bitmap <= 16'b0000000000000000;
		15'h0d0d: char_row_bitmap <= 16'b0000000000000000;
		15'h0d0e: char_row_bitmap <= 16'b0000000000000000;
		15'h0d0f: char_row_bitmap <= 16'b0000000000000000;
		15'h0d10: char_row_bitmap <= 16'b0000000000000000;
		15'h0d11: char_row_bitmap <= 16'b0001111000011000;
		15'h0d12: char_row_bitmap <= 16'b0011111100111000;
		15'h0d13: char_row_bitmap <= 16'b0111001111110000;
		15'h0d14: char_row_bitmap <= 16'b0110001111100000;
		15'h0d15: char_row_bitmap <= 16'b0000001100000000;
		15'h0d16: char_row_bitmap <= 16'b0000001100000000;
		15'h0d17: char_row_bitmap <= 16'b0000001100000000;
		15'h0d18: char_row_bitmap <= 16'b0000001100000000;
		15'h0d19: char_row_bitmap <= 16'b0000001100000000;
		15'h0d1a: char_row_bitmap <= 16'b0000001100000000;
		15'h0d1b: char_row_bitmap <= 16'b0000001100000000;
		15'h0d1c: char_row_bitmap <= 16'b0000000000000000;
		15'h0d1d: char_row_bitmap <= 16'b0000000000000000;
		15'h0d1e: char_row_bitmap <= 16'b0000000000000000;
		15'h0d1f: char_row_bitmap <= 16'b0000000000000000;
		15'h0d20: char_row_bitmap <= 16'b0000000000000000;
		15'h0d21: char_row_bitmap <= 16'b0000000000000000;
		15'h0d22: char_row_bitmap <= 16'b0000011110000000;
		15'h0d23: char_row_bitmap <= 16'b0000111111000000;
		15'h0d24: char_row_bitmap <= 16'b0001110011100000;
		15'h0d25: char_row_bitmap <= 16'b0001100001100000;
		15'h0d26: char_row_bitmap <= 16'b0011000000110000;
		15'h0d27: char_row_bitmap <= 16'b0011000000110000;
		15'h0d28: char_row_bitmap <= 16'b0011111111110000;
		15'h0d29: char_row_bitmap <= 16'b0011111111110000;
		15'h0d2a: char_row_bitmap <= 16'b0011000000110000;
		15'h0d2b: char_row_bitmap <= 16'b0011000000110000;
		15'h0d2c: char_row_bitmap <= 16'b0001100001100000;
		15'h0d2d: char_row_bitmap <= 16'b0001110011100000;
		15'h0d2e: char_row_bitmap <= 16'b0000111111000000;
		15'h0d2f: char_row_bitmap <= 16'b0000011110000000;
		15'h0d30: char_row_bitmap <= 16'b0000000000000000;
		15'h0d31: char_row_bitmap <= 16'b0000000000000000;
		15'h0d32: char_row_bitmap <= 16'b0000000000000000;
		15'h0d33: char_row_bitmap <= 16'b0000000000000000;
		15'h0d34: char_row_bitmap <= 16'b0000000000000000;
		15'h0d35: char_row_bitmap <= 16'b0000000000000000;
		15'h0d36: char_row_bitmap <= 16'b0000000000000000;
		15'h0d37: char_row_bitmap <= 16'b0000111111000000;
		15'h0d38: char_row_bitmap <= 16'b0001111111100000;
		15'h0d39: char_row_bitmap <= 16'b0011100001110000;
		15'h0d3a: char_row_bitmap <= 16'b0011000000110000;
		15'h0d3b: char_row_bitmap <= 16'b0011000000110000;
		15'h0d3c: char_row_bitmap <= 16'b0011000000110000;
		15'h0d3d: char_row_bitmap <= 16'b0011000000110000;
		15'h0d3e: char_row_bitmap <= 16'b0011100001110000;
		15'h0d3f: char_row_bitmap <= 16'b0001110011100000;
		15'h0d40: char_row_bitmap <= 16'b0000110011000000;
		15'h0d41: char_row_bitmap <= 16'b0000110011000000;
		15'h0d42: char_row_bitmap <= 16'b0011110011110000;
		15'h0d43: char_row_bitmap <= 16'b0011110011110000;
		15'h0d44: char_row_bitmap <= 16'b0000000000000000;
		15'h0d45: char_row_bitmap <= 16'b0000000000000000;
		15'h0d46: char_row_bitmap <= 16'b0000000000000000;
		15'h0d47: char_row_bitmap <= 16'b0000000000000000;
		15'h0d48: char_row_bitmap <= 16'b0000000000000000;
		15'h0d49: char_row_bitmap <= 16'b0000000000000000;
		15'h0d4a: char_row_bitmap <= 16'b0000000001100000;
		15'h0d4b: char_row_bitmap <= 16'b0000000111100000;
		15'h0d4c: char_row_bitmap <= 16'b0000001111000000;
		15'h0d4d: char_row_bitmap <= 16'b0000001100000000;
		15'h0d4e: char_row_bitmap <= 16'b0000001100000000;
		15'h0d4f: char_row_bitmap <= 16'b0000001110000000;
		15'h0d50: char_row_bitmap <= 16'b0000111110000000;
		15'h0d51: char_row_bitmap <= 16'b0001111111000000;
		15'h0d52: char_row_bitmap <= 16'b0011100111000000;
		15'h0d53: char_row_bitmap <= 16'b0011000011000000;
		15'h0d54: char_row_bitmap <= 16'b0011000011000000;
		15'h0d55: char_row_bitmap <= 16'b0011100111000000;
		15'h0d56: char_row_bitmap <= 16'b0001111110000000;
		15'h0d57: char_row_bitmap <= 16'b0000111100000000;
		15'h0d58: char_row_bitmap <= 16'b0000000000000000;
		15'h0d59: char_row_bitmap <= 16'b0000000000000000;
		15'h0d5a: char_row_bitmap <= 16'b0000000000000000;
		15'h0d5b: char_row_bitmap <= 16'b0000000000000000;
		15'h0d5c: char_row_bitmap <= 16'b0000000000000000;
		15'h0d5d: char_row_bitmap <= 16'b0000000000000000;
		15'h0d5e: char_row_bitmap <= 16'b0000000000000000;
		15'h0d5f: char_row_bitmap <= 16'b0000000000000000;
		15'h0d60: char_row_bitmap <= 16'b0000000100000000;
		15'h0d61: char_row_bitmap <= 16'b0000000100000000;
		15'h0d62: char_row_bitmap <= 16'b0000001110000000;
		15'h0d63: char_row_bitmap <= 16'b0000001110000000;
		15'h0d64: char_row_bitmap <= 16'b0000011011000000;
		15'h0d65: char_row_bitmap <= 16'b0000011011000000;
		15'h0d66: char_row_bitmap <= 16'b0000110001100000;
		15'h0d67: char_row_bitmap <= 16'b0000110001100000;
		15'h0d68: char_row_bitmap <= 16'b0001100000110000;
		15'h0d69: char_row_bitmap <= 16'b0001100000110000;
		15'h0d6a: char_row_bitmap <= 16'b0011111111111000;
		15'h0d6b: char_row_bitmap <= 16'b0011111111111000;
		15'h0d6c: char_row_bitmap <= 16'b0000000000000000;
		15'h0d6d: char_row_bitmap <= 16'b0000000000000000;
		15'h0d6e: char_row_bitmap <= 16'b0000000000000000;
		15'h0d6f: char_row_bitmap <= 16'b0000000000000000;
		15'h0d70: char_row_bitmap <= 16'b0000000000000000;
		15'h0d71: char_row_bitmap <= 16'b0000000000000000;
		15'h0d72: char_row_bitmap <= 16'b0000000000000000;
		15'h0d73: char_row_bitmap <= 16'b0000000000000000;
		15'h0d74: char_row_bitmap <= 16'b0000000000000000;
		15'h0d75: char_row_bitmap <= 16'b0000000000000000;
		15'h0d76: char_row_bitmap <= 16'b0000111111000000;
		15'h0d77: char_row_bitmap <= 16'b0001111111000000;
		15'h0d78: char_row_bitmap <= 16'b0011100000000000;
		15'h0d79: char_row_bitmap <= 16'b0011000000000000;
		15'h0d7a: char_row_bitmap <= 16'b0011111111000000;
		15'h0d7b: char_row_bitmap <= 16'b0011111111000000;
		15'h0d7c: char_row_bitmap <= 16'b0011000000000000;
		15'h0d7d: char_row_bitmap <= 16'b0011100000000000;
		15'h0d7e: char_row_bitmap <= 16'b0001111111000000;
		15'h0d7f: char_row_bitmap <= 16'b0000111111000000;
		15'h0d80: char_row_bitmap <= 16'b0000000000000000;
		15'h0d81: char_row_bitmap <= 16'b0000000000000000;
		15'h0d82: char_row_bitmap <= 16'b0000000000000000;
		15'h0d83: char_row_bitmap <= 16'b0000000000000000;
		15'h0d84: char_row_bitmap <= 16'b0000000000000000;
		15'h0d85: char_row_bitmap <= 16'b0000000000000000;
		15'h0d86: char_row_bitmap <= 16'b0000000000000000;
		15'h0d87: char_row_bitmap <= 16'b0011000001100000;
		15'h0d88: char_row_bitmap <= 16'b0011000001100000;
		15'h0d89: char_row_bitmap <= 16'b0011000001100000;
		15'h0d8a: char_row_bitmap <= 16'b0011000001100000;
		15'h0d8b: char_row_bitmap <= 16'b0011000001100000;
		15'h0d8c: char_row_bitmap <= 16'b0011000001100000;
		15'h0d8d: char_row_bitmap <= 16'b0011000001100000;
		15'h0d8e: char_row_bitmap <= 16'b0011000001100000;
		15'h0d8f: char_row_bitmap <= 16'b0011000001100000;
		15'h0d90: char_row_bitmap <= 16'b0011000001100000;
		15'h0d91: char_row_bitmap <= 16'b0011100011100000;
		15'h0d92: char_row_bitmap <= 16'b0001111111000000;
		15'h0d93: char_row_bitmap <= 16'b0000111110000000;
		15'h0d94: char_row_bitmap <= 16'b0000000000000000;
		15'h0d95: char_row_bitmap <= 16'b0000000000000000;
		15'h0d96: char_row_bitmap <= 16'b0000000000000000;
		15'h0d97: char_row_bitmap <= 16'b0000000000000000;
		15'h0d98: char_row_bitmap <= 16'b0000000000000000;
		15'h0d99: char_row_bitmap <= 16'b0000000000000000;
		15'h0d9a: char_row_bitmap <= 16'b0000000000000000;
		15'h0d9b: char_row_bitmap <= 16'b0000111110000000;
		15'h0d9c: char_row_bitmap <= 16'b0001111111000000;
		15'h0d9d: char_row_bitmap <= 16'b0011100011100000;
		15'h0d9e: char_row_bitmap <= 16'b0011000001100000;
		15'h0d9f: char_row_bitmap <= 16'b0011000001100000;
		15'h0da0: char_row_bitmap <= 16'b0011000001100000;
		15'h0da1: char_row_bitmap <= 16'b0011000001100000;
		15'h0da2: char_row_bitmap <= 16'b0011000001100000;
		15'h0da3: char_row_bitmap <= 16'b0011000001100000;
		15'h0da4: char_row_bitmap <= 16'b0011000001100000;
		15'h0da5: char_row_bitmap <= 16'b0011000001100000;
		15'h0da6: char_row_bitmap <= 16'b0011000001100000;
		15'h0da7: char_row_bitmap <= 16'b0011000001100000;
		15'h0da8: char_row_bitmap <= 16'b0000000000000000;
		15'h0da9: char_row_bitmap <= 16'b0000000000000000;
		15'h0daa: char_row_bitmap <= 16'b0000000000000000;
		15'h0dab: char_row_bitmap <= 16'b0000000000000000;
		15'h0dac: char_row_bitmap <= 16'b0000000000000000;
		15'h0dad: char_row_bitmap <= 16'b0000000000000000;
		15'h0dae: char_row_bitmap <= 16'b0000000000000000;
		15'h0daf: char_row_bitmap <= 16'b0000000000000000;
		15'h0db0: char_row_bitmap <= 16'b0000000000000000;
		15'h0db1: char_row_bitmap <= 16'b0000000000000000;
		15'h0db2: char_row_bitmap <= 16'b0000000000000000;
		15'h0db3: char_row_bitmap <= 16'b0000111001110000;
		15'h0db4: char_row_bitmap <= 16'b0001111111111000;
		15'h0db5: char_row_bitmap <= 16'b0011101110011100;
		15'h0db6: char_row_bitmap <= 16'b0011000110001100;
		15'h0db7: char_row_bitmap <= 16'b0011000110001100;
		15'h0db8: char_row_bitmap <= 16'b0011000110001100;
		15'h0db9: char_row_bitmap <= 16'b0011101111011100;
		15'h0dba: char_row_bitmap <= 16'b0001111111111000;
		15'h0dbb: char_row_bitmap <= 16'b0000111001110000;
		15'h0dbc: char_row_bitmap <= 16'b0000000000000000;
		15'h0dbd: char_row_bitmap <= 16'b0000000000000000;
		15'h0dbe: char_row_bitmap <= 16'b0000000000000000;
		15'h0dbf: char_row_bitmap <= 16'b0000000000000000;
		15'h0dc0: char_row_bitmap <= 16'b0000000000000000;
		15'h0dc1: char_row_bitmap <= 16'b0000000000000000;
		15'h0dc2: char_row_bitmap <= 16'b0000000110000000;
		15'h0dc3: char_row_bitmap <= 16'b0000001111000000;
		15'h0dc4: char_row_bitmap <= 16'b0000011111100000;
		15'h0dc5: char_row_bitmap <= 16'b0000011001100000;
		15'h0dc6: char_row_bitmap <= 16'b0000011001100000;
		15'h0dc7: char_row_bitmap <= 16'b0000011111100000;
		15'h0dc8: char_row_bitmap <= 16'b0000001111000000;
		15'h0dc9: char_row_bitmap <= 16'b0000000110000000;
		15'h0dca: char_row_bitmap <= 16'b0000000000000000;
		15'h0dcb: char_row_bitmap <= 16'b0000000000000000;
		15'h0dcc: char_row_bitmap <= 16'b0000000000000000;
		15'h0dcd: char_row_bitmap <= 16'b0000000000000000;
		15'h0dce: char_row_bitmap <= 16'b0000000000000000;
		15'h0dcf: char_row_bitmap <= 16'b0000000000000000;
		15'h0dd0: char_row_bitmap <= 16'b0000000000000000;
		15'h0dd1: char_row_bitmap <= 16'b0000000000000000;
		15'h0dd2: char_row_bitmap <= 16'b0000000000000000;
		15'h0dd3: char_row_bitmap <= 16'b0000000000000000;
		15'h0dd4: char_row_bitmap <= 16'b0000000000000000;
		15'h0dd5: char_row_bitmap <= 16'b0000000000000000;
		15'h0dd6: char_row_bitmap <= 16'b0000000110000000;
		15'h0dd7: char_row_bitmap <= 16'b0000001110000000;
		15'h0dd8: char_row_bitmap <= 16'b0000011110000000;
		15'h0dd9: char_row_bitmap <= 16'b0000000110000000;
		15'h0dda: char_row_bitmap <= 16'b0000000110000000;
		15'h0ddb: char_row_bitmap <= 16'b0000000110000000;
		15'h0ddc: char_row_bitmap <= 16'b0000000110000000;
		15'h0ddd: char_row_bitmap <= 16'b0000000110000000;
		15'h0dde: char_row_bitmap <= 16'b0000000000000000;
		15'h0ddf: char_row_bitmap <= 16'b0000000000000000;
		15'h0de0: char_row_bitmap <= 16'b0000000000000000;
		15'h0de1: char_row_bitmap <= 16'b0000000000000000;
		15'h0de2: char_row_bitmap <= 16'b0000000000000000;
		15'h0de3: char_row_bitmap <= 16'b0000000000000000;
		15'h0de4: char_row_bitmap <= 16'b0000000000000000;
		15'h0de5: char_row_bitmap <= 16'b0000000000000000;
		15'h0de6: char_row_bitmap <= 16'b0000000000000000;
		15'h0de7: char_row_bitmap <= 16'b0000000000000000;
		15'h0de8: char_row_bitmap <= 16'b0000000000000000;
		15'h0de9: char_row_bitmap <= 16'b0000000000000000;
		15'h0dea: char_row_bitmap <= 16'b0000011111100000;
		15'h0deb: char_row_bitmap <= 16'b0000111111110000;
		15'h0dec: char_row_bitmap <= 16'b0000110001110000;
		15'h0ded: char_row_bitmap <= 16'b0000000111100000;
		15'h0dee: char_row_bitmap <= 16'b0000001111000000;
		15'h0def: char_row_bitmap <= 16'b0000011100000000;
		15'h0df0: char_row_bitmap <= 16'b0000111111110000;
		15'h0df1: char_row_bitmap <= 16'b0000111111110000;
		15'h0df2: char_row_bitmap <= 16'b0000000000000000;
		15'h0df3: char_row_bitmap <= 16'b0000000000000000;
		15'h0df4: char_row_bitmap <= 16'b0000000000000000;
		15'h0df5: char_row_bitmap <= 16'b0000000000000000;
		15'h0df6: char_row_bitmap <= 16'b0000000000000000;
		15'h0df7: char_row_bitmap <= 16'b0000000000000000;
		15'h0df8: char_row_bitmap <= 16'b0000000000000000;
		15'h0df9: char_row_bitmap <= 16'b0000000000000000;
		15'h0dfa: char_row_bitmap <= 16'b0000000000000000;
		15'h0dfb: char_row_bitmap <= 16'b0000000000000000;
		15'h0dfc: char_row_bitmap <= 16'b0000000000000000;
		15'h0dfd: char_row_bitmap <= 16'b0000000000000000;
		15'h0dfe: char_row_bitmap <= 16'b0000011111100000;
		15'h0dff: char_row_bitmap <= 16'b0000011111110000;
		15'h0e00: char_row_bitmap <= 16'b0000000001110000;
		15'h0e01: char_row_bitmap <= 16'b0000000111100000;
		15'h0e02: char_row_bitmap <= 16'b0000000111100000;
		15'h0e03: char_row_bitmap <= 16'b0000000001110000;
		15'h0e04: char_row_bitmap <= 16'b0000011111110000;
		15'h0e05: char_row_bitmap <= 16'b0000011111100000;
		15'h0e06: char_row_bitmap <= 16'b0000000000000000;
		15'h0e07: char_row_bitmap <= 16'b0000000000000000;
		15'h0e08: char_row_bitmap <= 16'b0000000000000000;
		15'h0e09: char_row_bitmap <= 16'b0000000000000000;
		15'h0e0a: char_row_bitmap <= 16'b0000000000000000;
		15'h0e0b: char_row_bitmap <= 16'b0000000000000000;
		15'h0e0c: char_row_bitmap <= 16'b0000000000000000;
		15'h0e0d: char_row_bitmap <= 16'b0000000000000000;
		15'h0e0e: char_row_bitmap <= 16'b0000000000000000;
		15'h0e0f: char_row_bitmap <= 16'b0000000000000000;
		15'h0e10: char_row_bitmap <= 16'b0000000000000000;
		15'h0e11: char_row_bitmap <= 16'b0000000000000000;
		15'h0e12: char_row_bitmap <= 16'b0000000011000000;
		15'h0e13: char_row_bitmap <= 16'b0000000111000000;
		15'h0e14: char_row_bitmap <= 16'b0000001111000000;
		15'h0e15: char_row_bitmap <= 16'b0000011011000000;
		15'h0e16: char_row_bitmap <= 16'b0000111111110000;
		15'h0e17: char_row_bitmap <= 16'b0000111111110000;
		15'h0e18: char_row_bitmap <= 16'b0000000011000000;
		15'h0e19: char_row_bitmap <= 16'b0000000011000000;
		15'h0e1a: char_row_bitmap <= 16'b0000000000000000;
		15'h0e1b: char_row_bitmap <= 16'b0000000000000000;
		15'h0e1c: char_row_bitmap <= 16'b0000000000000000;
		15'h0e1d: char_row_bitmap <= 16'b0000000000000000;
		15'h0e1e: char_row_bitmap <= 16'b0000000000000000;
		15'h0e1f: char_row_bitmap <= 16'b0000000000000000;
		15'h0e20: char_row_bitmap <= 16'b0000000000000000;
		15'h0e21: char_row_bitmap <= 16'b0000000000000000;
		15'h0e22: char_row_bitmap <= 16'b0000000000000000;
		15'h0e23: char_row_bitmap <= 16'b0000000000000000;
		15'h0e24: char_row_bitmap <= 16'b0000000000000000;
		15'h0e25: char_row_bitmap <= 16'b0000000000000000;
		15'h0e26: char_row_bitmap <= 16'b0000111111110000;
		15'h0e27: char_row_bitmap <= 16'b0000111111110000;
		15'h0e28: char_row_bitmap <= 16'b0000110000000000;
		15'h0e29: char_row_bitmap <= 16'b0000111111100000;
		15'h0e2a: char_row_bitmap <= 16'b0000111111110000;
		15'h0e2b: char_row_bitmap <= 16'b0000000000110000;
		15'h0e2c: char_row_bitmap <= 16'b0000111111110000;
		15'h0e2d: char_row_bitmap <= 16'b0000011111100000;
		15'h0e2e: char_row_bitmap <= 16'b0000000000000000;
		15'h0e2f: char_row_bitmap <= 16'b0000000000000000;
		15'h0e30: char_row_bitmap <= 16'b0000000000000000;
		15'h0e31: char_row_bitmap <= 16'b0000000000000000;
		15'h0e32: char_row_bitmap <= 16'b0000000000000000;
		15'h0e33: char_row_bitmap <= 16'b0000000000000000;
		15'h0e34: char_row_bitmap <= 16'b0000000000000000;
		15'h0e35: char_row_bitmap <= 16'b0000000000000000;
		15'h0e36: char_row_bitmap <= 16'b0000000000000000;
		15'h0e37: char_row_bitmap <= 16'b0000000000000000;
		15'h0e38: char_row_bitmap <= 16'b0000000000000000;
		15'h0e39: char_row_bitmap <= 16'b0000000000000000;
		15'h0e3a: char_row_bitmap <= 16'b0000001111100000;
		15'h0e3b: char_row_bitmap <= 16'b0000011111100000;
		15'h0e3c: char_row_bitmap <= 16'b0000111000000000;
		15'h0e3d: char_row_bitmap <= 16'b0000111111100000;
		15'h0e3e: char_row_bitmap <= 16'b0000111111110000;
		15'h0e3f: char_row_bitmap <= 16'b0000110000110000;
		15'h0e40: char_row_bitmap <= 16'b0000111111110000;
		15'h0e41: char_row_bitmap <= 16'b0000011111100000;
		15'h0e42: char_row_bitmap <= 16'b0000000000000000;
		15'h0e43: char_row_bitmap <= 16'b0000000000000000;
		15'h0e44: char_row_bitmap <= 16'b0000000000000000;
		15'h0e45: char_row_bitmap <= 16'b0000000000000000;
		15'h0e46: char_row_bitmap <= 16'b0000000000000000;
		15'h0e47: char_row_bitmap <= 16'b0000000000000000;
		15'h0e48: char_row_bitmap <= 16'b0000000000000000;
		15'h0e49: char_row_bitmap <= 16'b0000000000000000;
		15'h0e4a: char_row_bitmap <= 16'b0000000000000000;
		15'h0e4b: char_row_bitmap <= 16'b0000000000000000;
		15'h0e4c: char_row_bitmap <= 16'b0000000000000000;
		15'h0e4d: char_row_bitmap <= 16'b0000000000000000;
		15'h0e4e: char_row_bitmap <= 16'b0000111111110000;
		15'h0e4f: char_row_bitmap <= 16'b0000111111110000;
		15'h0e50: char_row_bitmap <= 16'b0000000001110000;
		15'h0e51: char_row_bitmap <= 16'b0000000011100000;
		15'h0e52: char_row_bitmap <= 16'b0000000111000000;
		15'h0e53: char_row_bitmap <= 16'b0000000110000000;
		15'h0e54: char_row_bitmap <= 16'b0000000110000000;
		15'h0e55: char_row_bitmap <= 16'b0000000110000000;
		15'h0e56: char_row_bitmap <= 16'b0000000000000000;
		15'h0e57: char_row_bitmap <= 16'b0000000000000000;
		15'h0e58: char_row_bitmap <= 16'b0000000000000000;
		15'h0e59: char_row_bitmap <= 16'b0000000000000000;
		15'h0e5a: char_row_bitmap <= 16'b0000000000000000;
		15'h0e5b: char_row_bitmap <= 16'b0000000000000000;
		15'h0e5c: char_row_bitmap <= 16'b0000000000000000;
		15'h0e5d: char_row_bitmap <= 16'b0000000000000000;
		15'h0e5e: char_row_bitmap <= 16'b0000000000000000;
		15'h0e5f: char_row_bitmap <= 16'b0000000000000000;
		15'h0e60: char_row_bitmap <= 16'b0000000000000000;
		15'h0e61: char_row_bitmap <= 16'b0000000000000000;
		15'h0e62: char_row_bitmap <= 16'b0000011111100000;
		15'h0e63: char_row_bitmap <= 16'b0000111111110000;
		15'h0e64: char_row_bitmap <= 16'b0000110000110000;
		15'h0e65: char_row_bitmap <= 16'b0000011111100000;
		15'h0e66: char_row_bitmap <= 16'b0000111111110000;
		15'h0e67: char_row_bitmap <= 16'b0000110000110000;
		15'h0e68: char_row_bitmap <= 16'b0000111111110000;
		15'h0e69: char_row_bitmap <= 16'b0000011111100000;
		15'h0e6a: char_row_bitmap <= 16'b0000000000000000;
		15'h0e6b: char_row_bitmap <= 16'b0000000000000000;
		15'h0e6c: char_row_bitmap <= 16'b0000000000000000;
		15'h0e6d: char_row_bitmap <= 16'b0000000000000000;
		15'h0e6e: char_row_bitmap <= 16'b0000000000000000;
		15'h0e6f: char_row_bitmap <= 16'b0000000000000000;
		15'h0e70: char_row_bitmap <= 16'b0000000000000000;
		15'h0e71: char_row_bitmap <= 16'b0000000000000000;
		15'h0e72: char_row_bitmap <= 16'b0000000000000000;
		15'h0e73: char_row_bitmap <= 16'b0000000000000000;
		15'h0e74: char_row_bitmap <= 16'b0000000000000000;
		15'h0e75: char_row_bitmap <= 16'b0000000000000000;
		15'h0e76: char_row_bitmap <= 16'b0000011111100000;
		15'h0e77: char_row_bitmap <= 16'b0000111111110000;
		15'h0e78: char_row_bitmap <= 16'b0000110000110000;
		15'h0e79: char_row_bitmap <= 16'b0000111111110000;
		15'h0e7a: char_row_bitmap <= 16'b0000011111110000;
		15'h0e7b: char_row_bitmap <= 16'b0000000000110000;
		15'h0e7c: char_row_bitmap <= 16'b0000011111110000;
		15'h0e7d: char_row_bitmap <= 16'b0000011111100000;
		15'h0e7e: char_row_bitmap <= 16'b0000000000000000;
		15'h0e7f: char_row_bitmap <= 16'b0000000000000000;
		15'h0e80: char_row_bitmap <= 16'b0000000000000000;
		15'h0e81: char_row_bitmap <= 16'b0000000000000000;
		15'h0e82: char_row_bitmap <= 16'b0000000000000000;
		15'h0e83: char_row_bitmap <= 16'b0000000000000000;
		15'h0e84: char_row_bitmap <= 16'b0000000000000000;
		15'h0e85: char_row_bitmap <= 16'b0000000000000000;
		15'h0e86: char_row_bitmap <= 16'b0000000000000000;
		15'h0e87: char_row_bitmap <= 16'b0000000000000000;
		15'h0e88: char_row_bitmap <= 16'b0000000000000000;
		15'h0e89: char_row_bitmap <= 16'b0000000000000000;
		15'h0e8a: char_row_bitmap <= 16'b0000000000110000;
		15'h0e8b: char_row_bitmap <= 16'b0000000001110000;
		15'h0e8c: char_row_bitmap <= 16'b0000000011100000;
		15'h0e8d: char_row_bitmap <= 16'b0000000111000000;
		15'h0e8e: char_row_bitmap <= 16'b0000001110000000;
		15'h0e8f: char_row_bitmap <= 16'b0000011100000000;
		15'h0e90: char_row_bitmap <= 16'b0000111000000000;
		15'h0e91: char_row_bitmap <= 16'b0001110000000000;
		15'h0e92: char_row_bitmap <= 16'b0000111000000000;
		15'h0e93: char_row_bitmap <= 16'b0000011100000000;
		15'h0e94: char_row_bitmap <= 16'b0011001110000000;
		15'h0e95: char_row_bitmap <= 16'b0011100111000000;
		15'h0e96: char_row_bitmap <= 16'b0001110011100000;
		15'h0e97: char_row_bitmap <= 16'b0000111001110000;
		15'h0e98: char_row_bitmap <= 16'b0000011100110000;
		15'h0e99: char_row_bitmap <= 16'b0000001110000000;
		15'h0e9a: char_row_bitmap <= 16'b0000000111000000;
		15'h0e9b: char_row_bitmap <= 16'b0000000011000000;
		15'h0e9c: char_row_bitmap <= 16'b0000000000000000;
		15'h0e9d: char_row_bitmap <= 16'b0000000000000000;
		15'h0e9e: char_row_bitmap <= 16'b0000000000000000;
		15'h0e9f: char_row_bitmap <= 16'b0000000000000000;
		15'h0ea0: char_row_bitmap <= 16'b0001111000011000;
		15'h0ea1: char_row_bitmap <= 16'b0011111100111000;
		15'h0ea2: char_row_bitmap <= 16'b0111001111110000;
		15'h0ea3: char_row_bitmap <= 16'b0110000111100000;
		15'h0ea4: char_row_bitmap <= 16'b0000000000000000;
		15'h0ea5: char_row_bitmap <= 16'b0000000000000000;
		15'h0ea6: char_row_bitmap <= 16'b0011111111110000;
		15'h0ea7: char_row_bitmap <= 16'b0011111111110000;
		15'h0ea8: char_row_bitmap <= 16'b0000000000000000;
		15'h0ea9: char_row_bitmap <= 16'b0000000000000000;
		15'h0eaa: char_row_bitmap <= 16'b0000000000000000;
		15'h0eab: char_row_bitmap <= 16'b0000000000000000;
		15'h0eac: char_row_bitmap <= 16'b0000000000000000;
		15'h0ead: char_row_bitmap <= 16'b0000000000000000;
		15'h0eae: char_row_bitmap <= 16'b0000000000000000;
		15'h0eaf: char_row_bitmap <= 16'b0000000000000000;
		15'h0eb0: char_row_bitmap <= 16'b0000000000000000;
		15'h0eb1: char_row_bitmap <= 16'b0000000000000000;
		15'h0eb2: char_row_bitmap <= 16'b0011000000000000;
		15'h0eb3: char_row_bitmap <= 16'b0011100000000000;
		15'h0eb4: char_row_bitmap <= 16'b0001110000000000;
		15'h0eb5: char_row_bitmap <= 16'b0000111000000000;
		15'h0eb6: char_row_bitmap <= 16'b0000011100000000;
		15'h0eb7: char_row_bitmap <= 16'b0000001110000000;
		15'h0eb8: char_row_bitmap <= 16'b0000000111000000;
		15'h0eb9: char_row_bitmap <= 16'b0000000011100000;
		15'h0eba: char_row_bitmap <= 16'b0000000111000000;
		15'h0ebb: char_row_bitmap <= 16'b0000001110000000;
		15'h0ebc: char_row_bitmap <= 16'b0000011100110000;
		15'h0ebd: char_row_bitmap <= 16'b0000111001110000;
		15'h0ebe: char_row_bitmap <= 16'b0001110011100000;
		15'h0ebf: char_row_bitmap <= 16'b0011100111000000;
		15'h0ec0: char_row_bitmap <= 16'b0011001110000000;
		15'h0ec1: char_row_bitmap <= 16'b0000011100000000;
		15'h0ec2: char_row_bitmap <= 16'b0000111000000000;
		15'h0ec3: char_row_bitmap <= 16'b0000110000000000;
		15'h0ec4: char_row_bitmap <= 16'b0000000000000000;
		15'h0ec5: char_row_bitmap <= 16'b0000000000000000;
		15'h0ec6: char_row_bitmap <= 16'b0000000000000000;
		15'h0ec7: char_row_bitmap <= 16'b0000000000000000;
		15'h0ec8: char_row_bitmap <= 16'b0000000000000000;
		15'h0ec9: char_row_bitmap <= 16'b0000000000000000;
		15'h0eca: char_row_bitmap <= 16'b0000000011001100;
		15'h0ecb: char_row_bitmap <= 16'b0000000111011100;
		15'h0ecc: char_row_bitmap <= 16'b0000001110111000;
		15'h0ecd: char_row_bitmap <= 16'b0000011101110000;
		15'h0ece: char_row_bitmap <= 16'b0000111011100000;
		15'h0ecf: char_row_bitmap <= 16'b0000011101110000;
		15'h0ed0: char_row_bitmap <= 16'b0000001110111000;
		15'h0ed1: char_row_bitmap <= 16'b0000000111011100;
		15'h0ed2: char_row_bitmap <= 16'b0000000011001100;
		15'h0ed3: char_row_bitmap <= 16'b0000000000000000;
		15'h0ed4: char_row_bitmap <= 16'b0000000000000000;
		15'h0ed5: char_row_bitmap <= 16'b0000000000000000;
		15'h0ed6: char_row_bitmap <= 16'b0000000000000000;
		15'h0ed7: char_row_bitmap <= 16'b0000000000000000;
		15'h0ed8: char_row_bitmap <= 16'b0000000000000000;
		15'h0ed9: char_row_bitmap <= 16'b0000000000000000;
		15'h0eda: char_row_bitmap <= 16'b0000000000000000;
		15'h0edb: char_row_bitmap <= 16'b0000000000000000;
		15'h0edc: char_row_bitmap <= 16'b0000000000000000;
		15'h0edd: char_row_bitmap <= 16'b0000000000000000;
		15'h0ede: char_row_bitmap <= 16'b0011001100000000;
		15'h0edf: char_row_bitmap <= 16'b0011101110000000;
		15'h0ee0: char_row_bitmap <= 16'b0001110111000000;
		15'h0ee1: char_row_bitmap <= 16'b0000111011100000;
		15'h0ee2: char_row_bitmap <= 16'b0000011101110000;
		15'h0ee3: char_row_bitmap <= 16'b0000111011100000;
		15'h0ee4: char_row_bitmap <= 16'b0001110111000000;
		15'h0ee5: char_row_bitmap <= 16'b0011101110000000;
		15'h0ee6: char_row_bitmap <= 16'b0011001100000000;
		15'h0ee7: char_row_bitmap <= 16'b0000000000000000;
		15'h0ee8: char_row_bitmap <= 16'b0000000000000000;
		15'h0ee9: char_row_bitmap <= 16'b0000000000000000;
		15'h0eea: char_row_bitmap <= 16'b0000000000000000;
		15'h0eeb: char_row_bitmap <= 16'b0000000000000000;
		15'h0eec: char_row_bitmap <= 16'b0000000000000000;
		15'h0eed: char_row_bitmap <= 16'b0000000000000000;
		15'h0eee: char_row_bitmap <= 16'b0001111111111100;
		15'h0eef: char_row_bitmap <= 16'b0011111111111100;
		15'h0ef0: char_row_bitmap <= 16'b0011000110110000;
		15'h0ef1: char_row_bitmap <= 16'b0011000110110000;
		15'h0ef2: char_row_bitmap <= 16'b0011000110110000;
		15'h0ef3: char_row_bitmap <= 16'b0011000110110000;
		15'h0ef4: char_row_bitmap <= 16'b0011111110110000;
		15'h0ef5: char_row_bitmap <= 16'b0001111110110000;
		15'h0ef6: char_row_bitmap <= 16'b0000000110110000;
		15'h0ef7: char_row_bitmap <= 16'b0000000110110000;
		15'h0ef8: char_row_bitmap <= 16'b0000000110110000;
		15'h0ef9: char_row_bitmap <= 16'b0000000110110000;
		15'h0efa: char_row_bitmap <= 16'b0000000110110000;
		15'h0efb: char_row_bitmap <= 16'b0000000110110000;
		15'h0efc: char_row_bitmap <= 16'b0000000110110000;
		15'h0efd: char_row_bitmap <= 16'b0000000000000000;
		15'h0efe: char_row_bitmap <= 16'b0000000000000000;
		15'h0eff: char_row_bitmap <= 16'b0000000000000000;
		15'h0f00: char_row_bitmap <= 16'b0000000000000000;
		15'h0f01: char_row_bitmap <= 16'b0000000000000000;
		15'h0f02: char_row_bitmap <= 16'b0000000000000000;
		15'h0f03: char_row_bitmap <= 16'b0000000000000000;
		15'h0f04: char_row_bitmap <= 16'b0000000000000000;
		15'h0f05: char_row_bitmap <= 16'b0000011100000000;
		15'h0f06: char_row_bitmap <= 16'b0000100000000000;
		15'h0f07: char_row_bitmap <= 16'b0000011000000000;
		15'h0f08: char_row_bitmap <= 16'b0000000100000000;
		15'h0f09: char_row_bitmap <= 16'b0000111000000000;
		15'h0f0a: char_row_bitmap <= 16'b0000000000000000;
		15'h0f0b: char_row_bitmap <= 16'b0000000001110000;
		15'h0f0c: char_row_bitmap <= 16'b0000000001001000;
		15'h0f0d: char_row_bitmap <= 16'b0000000001110000;
		15'h0f0e: char_row_bitmap <= 16'b0000000001000000;
		15'h0f0f: char_row_bitmap <= 16'b0000000001000000;
		15'h0f10: char_row_bitmap <= 16'b0000000000000000;
		15'h0f11: char_row_bitmap <= 16'b0000000000000000;
		15'h0f12: char_row_bitmap <= 16'b0000000000000000;
		15'h0f13: char_row_bitmap <= 16'b0000000000000000;
		15'h0f14: char_row_bitmap <= 16'b0000000000000000;
		15'h0f15: char_row_bitmap <= 16'b0000000000000000;
		15'h0f16: char_row_bitmap <= 16'b0000000000000000;
		15'h0f17: char_row_bitmap <= 16'b0000000000000000;
		15'h0f18: char_row_bitmap <= 16'b0000000000000000;
		15'h0f19: char_row_bitmap <= 16'b0000000000000000;
		15'h0f1a: char_row_bitmap <= 16'b0000111111000000;
		15'h0f1b: char_row_bitmap <= 16'b0001111111100000;
		15'h0f1c: char_row_bitmap <= 16'b0011100001110000;
		15'h0f1d: char_row_bitmap <= 16'b0011000000110000;
		15'h0f1e: char_row_bitmap <= 16'b0011111111110000;
		15'h0f1f: char_row_bitmap <= 16'b0011111111110000;
		15'h0f20: char_row_bitmap <= 16'b0011000000110000;
		15'h0f21: char_row_bitmap <= 16'b0011000000110000;
		15'h0f22: char_row_bitmap <= 16'b0011000000110000;
		15'h0f23: char_row_bitmap <= 16'b0011000000110000;
		15'h0f24: char_row_bitmap <= 16'b0000000000000000;
		15'h0f25: char_row_bitmap <= 16'b0000000000000000;
		15'h0f26: char_row_bitmap <= 16'b0000000000000000;
		15'h0f27: char_row_bitmap <= 16'b0000000000000000;
		15'h0f28: char_row_bitmap <= 16'b0000000000000000;
		15'h0f29: char_row_bitmap <= 16'b0000000000000000;
		15'h0f2a: char_row_bitmap <= 16'b0000000000000000;
		15'h0f2b: char_row_bitmap <= 16'b0000000000000000;
		15'h0f2c: char_row_bitmap <= 16'b0000000000000000;
		15'h0f2d: char_row_bitmap <= 16'b0000000000000000;
		15'h0f2e: char_row_bitmap <= 16'b0011111111000000;
		15'h0f2f: char_row_bitmap <= 16'b0011111111100000;
		15'h0f30: char_row_bitmap <= 16'b0011000001110000;
		15'h0f31: char_row_bitmap <= 16'b0011000001110000;
		15'h0f32: char_row_bitmap <= 16'b0011111111100000;
		15'h0f33: char_row_bitmap <= 16'b0011111111100000;
		15'h0f34: char_row_bitmap <= 16'b0011000001110000;
		15'h0f35: char_row_bitmap <= 16'b0011000001110000;
		15'h0f36: char_row_bitmap <= 16'b0011111111100000;
		15'h0f37: char_row_bitmap <= 16'b0011111111000000;
		15'h0f38: char_row_bitmap <= 16'b0000000000000000;
		15'h0f39: char_row_bitmap <= 16'b0000000000000000;
		15'h0f3a: char_row_bitmap <= 16'b0000000000000000;
		15'h0f3b: char_row_bitmap <= 16'b0000000000000000;
		15'h0f3c: char_row_bitmap <= 16'b0000000000000000;
		15'h0f3d: char_row_bitmap <= 16'b0000000000000000;
		15'h0f3e: char_row_bitmap <= 16'b0000000000000000;
		15'h0f3f: char_row_bitmap <= 16'b0000000000000000;
		15'h0f40: char_row_bitmap <= 16'b0000000000000000;
		15'h0f41: char_row_bitmap <= 16'b0000000000000000;
		15'h0f42: char_row_bitmap <= 16'b0000111111000000;
		15'h0f43: char_row_bitmap <= 16'b0001111111100000;
		15'h0f44: char_row_bitmap <= 16'b0011100001110000;
		15'h0f45: char_row_bitmap <= 16'b0011000000110000;
		15'h0f46: char_row_bitmap <= 16'b0011000000000000;
		15'h0f47: char_row_bitmap <= 16'b0011000000000000;
		15'h0f48: char_row_bitmap <= 16'b0011000000110000;
		15'h0f49: char_row_bitmap <= 16'b0011100001110000;
		15'h0f4a: char_row_bitmap <= 16'b0001111111100000;
		15'h0f4b: char_row_bitmap <= 16'b0000111111000000;
		15'h0f4c: char_row_bitmap <= 16'b0000000000000000;
		15'h0f4d: char_row_bitmap <= 16'b0000000000000000;
		15'h0f4e: char_row_bitmap <= 16'b0000000000000000;
		15'h0f4f: char_row_bitmap <= 16'b0000000000000000;
		15'h0f50: char_row_bitmap <= 16'b0000000000000000;
		15'h0f51: char_row_bitmap <= 16'b0000000000000000;
		15'h0f52: char_row_bitmap <= 16'b0000000000000000;
		15'h0f53: char_row_bitmap <= 16'b0000000000000000;
		15'h0f54: char_row_bitmap <= 16'b0000000000000000;
		15'h0f55: char_row_bitmap <= 16'b0000000000000000;
		15'h0f56: char_row_bitmap <= 16'b0011111111000000;
		15'h0f57: char_row_bitmap <= 16'b0011111111100000;
		15'h0f58: char_row_bitmap <= 16'b0011000001110000;
		15'h0f59: char_row_bitmap <= 16'b0011000000110000;
		15'h0f5a: char_row_bitmap <= 16'b0011000000110000;
		15'h0f5b: char_row_bitmap <= 16'b0011000000110000;
		15'h0f5c: char_row_bitmap <= 16'b0011000000110000;
		15'h0f5d: char_row_bitmap <= 16'b0011000001110000;
		15'h0f5e: char_row_bitmap <= 16'b0011111111100000;
		15'h0f5f: char_row_bitmap <= 16'b0011111111000000;
		15'h0f60: char_row_bitmap <= 16'b0000000000000000;
		15'h0f61: char_row_bitmap <= 16'b0000000000000000;
		15'h0f62: char_row_bitmap <= 16'b0000000000000000;
		15'h0f63: char_row_bitmap <= 16'b0000000000000000;
		15'h0f64: char_row_bitmap <= 16'b0000000000000000;
		15'h0f65: char_row_bitmap <= 16'b0000000000000000;
		15'h0f66: char_row_bitmap <= 16'b0000000000000000;
		15'h0f67: char_row_bitmap <= 16'b0000000000000000;
		15'h0f68: char_row_bitmap <= 16'b0000000000000000;
		15'h0f69: char_row_bitmap <= 16'b0000000000000000;
		15'h0f6a: char_row_bitmap <= 16'b0011111111110000;
		15'h0f6b: char_row_bitmap <= 16'b0011111111110000;
		15'h0f6c: char_row_bitmap <= 16'b0011000000000000;
		15'h0f6d: char_row_bitmap <= 16'b0011000000000000;
		15'h0f6e: char_row_bitmap <= 16'b0011111111000000;
		15'h0f6f: char_row_bitmap <= 16'b0011111111000000;
		15'h0f70: char_row_bitmap <= 16'b0011000000000000;
		15'h0f71: char_row_bitmap <= 16'b0011000000000000;
		15'h0f72: char_row_bitmap <= 16'b0011111111110000;
		15'h0f73: char_row_bitmap <= 16'b0011111111110000;
		15'h0f74: char_row_bitmap <= 16'b0000000000000000;
		15'h0f75: char_row_bitmap <= 16'b0000000000000000;
		15'h0f76: char_row_bitmap <= 16'b0000000000000000;
		15'h0f77: char_row_bitmap <= 16'b0000000000000000;
		15'h0f78: char_row_bitmap <= 16'b0000000000000000;
		15'h0f79: char_row_bitmap <= 16'b0000000000000000;
		15'h0f7a: char_row_bitmap <= 16'b0000000000000000;
		15'h0f7b: char_row_bitmap <= 16'b0000000000000000;
		15'h0f7c: char_row_bitmap <= 16'b0000000000000000;
		15'h0f7d: char_row_bitmap <= 16'b0000000000000000;
		15'h0f7e: char_row_bitmap <= 16'b0011111111110000;
		15'h0f7f: char_row_bitmap <= 16'b0011111111110000;
		15'h0f80: char_row_bitmap <= 16'b0011000000000000;
		15'h0f81: char_row_bitmap <= 16'b0011000000000000;
		15'h0f82: char_row_bitmap <= 16'b0011111111000000;
		15'h0f83: char_row_bitmap <= 16'b0011111111000000;
		15'h0f84: char_row_bitmap <= 16'b0011000000000000;
		15'h0f85: char_row_bitmap <= 16'b0011000000000000;
		15'h0f86: char_row_bitmap <= 16'b0011000000000000;
		15'h0f87: char_row_bitmap <= 16'b0011000000000000;
		15'h0f88: char_row_bitmap <= 16'b0000000000000000;
		15'h0f89: char_row_bitmap <= 16'b0000000000000000;
		15'h0f8a: char_row_bitmap <= 16'b0000000000000000;
		15'h0f8b: char_row_bitmap <= 16'b0000000000000000;
		15'h0f8c: char_row_bitmap <= 16'b0000000000000000;
		15'h0f8d: char_row_bitmap <= 16'b0000000000000000;
		15'h0f8e: char_row_bitmap <= 16'b0000000000000000;
		15'h0f8f: char_row_bitmap <= 16'b0000000000000000;
		15'h0f90: char_row_bitmap <= 16'b0000000000000000;
		15'h0f91: char_row_bitmap <= 16'b0000000000000000;
		15'h0f92: char_row_bitmap <= 16'b0000111111000000;
		15'h0f93: char_row_bitmap <= 16'b0001111111000000;
		15'h0f94: char_row_bitmap <= 16'b0011100000000000;
		15'h0f95: char_row_bitmap <= 16'b0011000000000000;
		15'h0f96: char_row_bitmap <= 16'b0011000011110000;
		15'h0f97: char_row_bitmap <= 16'b0011000011110000;
		15'h0f98: char_row_bitmap <= 16'b0011000000110000;
		15'h0f99: char_row_bitmap <= 16'b0011100000110000;
		15'h0f9a: char_row_bitmap <= 16'b0001111111110000;
		15'h0f9b: char_row_bitmap <= 16'b0000111111100000;
		15'h0f9c: char_row_bitmap <= 16'b0000000000000000;
		15'h0f9d: char_row_bitmap <= 16'b0000000000000000;
		15'h0f9e: char_row_bitmap <= 16'b0000000000000000;
		15'h0f9f: char_row_bitmap <= 16'b0000000000000000;
		15'h0fa0: char_row_bitmap <= 16'b0000000000000000;
		15'h0fa1: char_row_bitmap <= 16'b0000000000000000;
		15'h0fa2: char_row_bitmap <= 16'b0000000000000000;
		15'h0fa3: char_row_bitmap <= 16'b0000000000000000;
		15'h0fa4: char_row_bitmap <= 16'b0000000000000000;
		15'h0fa5: char_row_bitmap <= 16'b0000000000000000;
		15'h0fa6: char_row_bitmap <= 16'b0011000000110000;
		15'h0fa7: char_row_bitmap <= 16'b0011000000110000;
		15'h0fa8: char_row_bitmap <= 16'b0011000000110000;
		15'h0fa9: char_row_bitmap <= 16'b0011000000110000;
		15'h0faa: char_row_bitmap <= 16'b0011111111110000;
		15'h0fab: char_row_bitmap <= 16'b0011111111110000;
		15'h0fac: char_row_bitmap <= 16'b0011000000110000;
		15'h0fad: char_row_bitmap <= 16'b0011000000110000;
		15'h0fae: char_row_bitmap <= 16'b0011000000110000;
		15'h0faf: char_row_bitmap <= 16'b0011000000110000;
		15'h0fb0: char_row_bitmap <= 16'b0000000000000000;
		15'h0fb1: char_row_bitmap <= 16'b0000000000000000;
		15'h0fb2: char_row_bitmap <= 16'b0000000000000000;
		15'h0fb3: char_row_bitmap <= 16'b0000000000000000;
		15'h0fb4: char_row_bitmap <= 16'b0000000000000000;
		15'h0fb5: char_row_bitmap <= 16'b0000000000000000;
		15'h0fb6: char_row_bitmap <= 16'b0000000000000000;
		15'h0fb7: char_row_bitmap <= 16'b0000000000000000;
		15'h0fb8: char_row_bitmap <= 16'b0000000000000000;
		15'h0fb9: char_row_bitmap <= 16'b0000000000000000;
		15'h0fba: char_row_bitmap <= 16'b0000111111000000;
		15'h0fbb: char_row_bitmap <= 16'b0000111111000000;
		15'h0fbc: char_row_bitmap <= 16'b0000001100000000;
		15'h0fbd: char_row_bitmap <= 16'b0000001100000000;
		15'h0fbe: char_row_bitmap <= 16'b0000001100000000;
		15'h0fbf: char_row_bitmap <= 16'b0000001100000000;
		15'h0fc0: char_row_bitmap <= 16'b0000001100000000;
		15'h0fc1: char_row_bitmap <= 16'b0000001100000000;
		15'h0fc2: char_row_bitmap <= 16'b0000111111000000;
		15'h0fc3: char_row_bitmap <= 16'b0000111111000000;
		15'h0fc4: char_row_bitmap <= 16'b0000000000000000;
		15'h0fc5: char_row_bitmap <= 16'b0000000000000000;
		15'h0fc6: char_row_bitmap <= 16'b0000000000000000;
		15'h0fc7: char_row_bitmap <= 16'b0000000000000000;
		15'h0fc8: char_row_bitmap <= 16'b0000000000000000;
		15'h0fc9: char_row_bitmap <= 16'b0000000000000000;
		15'h0fca: char_row_bitmap <= 16'b0000000000000000;
		15'h0fcb: char_row_bitmap <= 16'b0000000000000000;
		15'h0fcc: char_row_bitmap <= 16'b0000000000000000;
		15'h0fcd: char_row_bitmap <= 16'b0000000000000000;
		15'h0fce: char_row_bitmap <= 16'b0000001111110000;
		15'h0fcf: char_row_bitmap <= 16'b0000001111110000;
		15'h0fd0: char_row_bitmap <= 16'b0000000011000000;
		15'h0fd1: char_row_bitmap <= 16'b0000000011000000;
		15'h0fd2: char_row_bitmap <= 16'b0000000011000000;
		15'h0fd3: char_row_bitmap <= 16'b0000000011000000;
		15'h0fd4: char_row_bitmap <= 16'b0011000011000000;
		15'h0fd5: char_row_bitmap <= 16'b0011100111000000;
		15'h0fd6: char_row_bitmap <= 16'b0001111110000000;
		15'h0fd7: char_row_bitmap <= 16'b0000111100000000;
		15'h0fd8: char_row_bitmap <= 16'b0000000000000000;
		15'h0fd9: char_row_bitmap <= 16'b0000000000000000;
		15'h0fda: char_row_bitmap <= 16'b0000000000000000;
		15'h0fdb: char_row_bitmap <= 16'b0000000000000000;
		15'h0fdc: char_row_bitmap <= 16'b0000000000000000;
		15'h0fdd: char_row_bitmap <= 16'b0000000000000000;
		15'h0fde: char_row_bitmap <= 16'b0000000000000000;
		15'h0fdf: char_row_bitmap <= 16'b0000000000000000;
		15'h0fe0: char_row_bitmap <= 16'b0000000000000000;
		15'h0fe1: char_row_bitmap <= 16'b0000000000000000;
		15'h0fe2: char_row_bitmap <= 16'b0011000000110000;
		15'h0fe3: char_row_bitmap <= 16'b0011000001110000;
		15'h0fe4: char_row_bitmap <= 16'b0011000011100000;
		15'h0fe5: char_row_bitmap <= 16'b0011000111000000;
		15'h0fe6: char_row_bitmap <= 16'b0011111110000000;
		15'h0fe7: char_row_bitmap <= 16'b0011111110000000;
		15'h0fe8: char_row_bitmap <= 16'b0011000111000000;
		15'h0fe9: char_row_bitmap <= 16'b0011000011100000;
		15'h0fea: char_row_bitmap <= 16'b0011000001110000;
		15'h0feb: char_row_bitmap <= 16'b0011000000110000;
		15'h0fec: char_row_bitmap <= 16'b0000000000000000;
		15'h0fed: char_row_bitmap <= 16'b0000000000000000;
		15'h0fee: char_row_bitmap <= 16'b0000000000000000;
		15'h0fef: char_row_bitmap <= 16'b0000000000000000;
		15'h0ff0: char_row_bitmap <= 16'b0000000000000000;
		15'h0ff1: char_row_bitmap <= 16'b0000000000000000;
		15'h0ff2: char_row_bitmap <= 16'b0000000000000000;
		15'h0ff3: char_row_bitmap <= 16'b0000000000000000;
		15'h0ff4: char_row_bitmap <= 16'b0000000000000000;
		15'h0ff5: char_row_bitmap <= 16'b0000000000000000;
		15'h0ff6: char_row_bitmap <= 16'b0011000000000000;
		15'h0ff7: char_row_bitmap <= 16'b0011000000000000;
		15'h0ff8: char_row_bitmap <= 16'b0011000000000000;
		15'h0ff9: char_row_bitmap <= 16'b0011000000000000;
		15'h0ffa: char_row_bitmap <= 16'b0011000000000000;
		15'h0ffb: char_row_bitmap <= 16'b0011000000000000;
		15'h0ffc: char_row_bitmap <= 16'b0011000000000000;
		15'h0ffd: char_row_bitmap <= 16'b0011000000000000;
		15'h0ffe: char_row_bitmap <= 16'b0011111111110000;
		15'h0fff: char_row_bitmap <= 16'b0011111111110000;
		15'h1000: char_row_bitmap <= 16'b0000000000000000;
		15'h1001: char_row_bitmap <= 16'b0000000000000000;
		15'h1002: char_row_bitmap <= 16'b0000000000000000;
		15'h1003: char_row_bitmap <= 16'b0000000000000000;
		15'h1004: char_row_bitmap <= 16'b0000000000000000;
		15'h1005: char_row_bitmap <= 16'b0000000000000000;
		15'h1006: char_row_bitmap <= 16'b0000000000000000;
		15'h1007: char_row_bitmap <= 16'b0000000000000000;
		15'h1008: char_row_bitmap <= 16'b0000000000000000;
		15'h1009: char_row_bitmap <= 16'b0000000000000000;
		15'h100a: char_row_bitmap <= 16'b0011000000110000;
		15'h100b: char_row_bitmap <= 16'b0011100001110000;
		15'h100c: char_row_bitmap <= 16'b0011110011110000;
		15'h100d: char_row_bitmap <= 16'b0011111111110000;
		15'h100e: char_row_bitmap <= 16'b0011011110110000;
		15'h100f: char_row_bitmap <= 16'b0011001100110000;
		15'h1010: char_row_bitmap <= 16'b0011000000110000;
		15'h1011: char_row_bitmap <= 16'b0011000000110000;
		15'h1012: char_row_bitmap <= 16'b0011000000110000;
		15'h1013: char_row_bitmap <= 16'b0011000000110000;
		15'h1014: char_row_bitmap <= 16'b0000000000000000;
		15'h1015: char_row_bitmap <= 16'b0000000000000000;
		15'h1016: char_row_bitmap <= 16'b0000000000000000;
		15'h1017: char_row_bitmap <= 16'b0000000000000000;
		15'h1018: char_row_bitmap <= 16'b0000000000000000;
		15'h1019: char_row_bitmap <= 16'b0000000000000000;
		15'h101a: char_row_bitmap <= 16'b0000000000000000;
		15'h101b: char_row_bitmap <= 16'b0000000000000000;
		15'h101c: char_row_bitmap <= 16'b0000000000000000;
		15'h101d: char_row_bitmap <= 16'b0000000000000000;
		15'h101e: char_row_bitmap <= 16'b0011000000110000;
		15'h101f: char_row_bitmap <= 16'b0011100000110000;
		15'h1020: char_row_bitmap <= 16'b0011110000110000;
		15'h1021: char_row_bitmap <= 16'b0011111000110000;
		15'h1022: char_row_bitmap <= 16'b0011011100110000;
		15'h1023: char_row_bitmap <= 16'b0011001110110000;
		15'h1024: char_row_bitmap <= 16'b0011000111110000;
		15'h1025: char_row_bitmap <= 16'b0011000011110000;
		15'h1026: char_row_bitmap <= 16'b0011000001110000;
		15'h1027: char_row_bitmap <= 16'b0011000000110000;
		15'h1028: char_row_bitmap <= 16'b0000000000000000;
		15'h1029: char_row_bitmap <= 16'b0000000000000000;
		15'h102a: char_row_bitmap <= 16'b0000000000000000;
		15'h102b: char_row_bitmap <= 16'b0000000000000000;
		15'h102c: char_row_bitmap <= 16'b0000000000000000;
		15'h102d: char_row_bitmap <= 16'b0000000000000000;
		15'h102e: char_row_bitmap <= 16'b0000000000000000;
		15'h102f: char_row_bitmap <= 16'b0000000000000000;
		15'h1030: char_row_bitmap <= 16'b0000000000000000;
		15'h1031: char_row_bitmap <= 16'b0000000000000000;
		15'h1032: char_row_bitmap <= 16'b0000111111000000;
		15'h1033: char_row_bitmap <= 16'b0001111111100000;
		15'h1034: char_row_bitmap <= 16'b0011100001110000;
		15'h1035: char_row_bitmap <= 16'b0011000000110000;
		15'h1036: char_row_bitmap <= 16'b0011000000110000;
		15'h1037: char_row_bitmap <= 16'b0011000000110000;
		15'h1038: char_row_bitmap <= 16'b0011000000110000;
		15'h1039: char_row_bitmap <= 16'b0011100001110000;
		15'h103a: char_row_bitmap <= 16'b0001111111100000;
		15'h103b: char_row_bitmap <= 16'b0000111111000000;
		15'h103c: char_row_bitmap <= 16'b0000000000000000;
		15'h103d: char_row_bitmap <= 16'b0000000000000000;
		15'h103e: char_row_bitmap <= 16'b0000000000000000;
		15'h103f: char_row_bitmap <= 16'b0000000000000000;
		15'h1040: char_row_bitmap <= 16'b0000000000000000;
		15'h1041: char_row_bitmap <= 16'b0000000000000000;
		15'h1042: char_row_bitmap <= 16'b0000000000000000;
		15'h1043: char_row_bitmap <= 16'b0000000000000000;
		15'h1044: char_row_bitmap <= 16'b0000000000000000;
		15'h1045: char_row_bitmap <= 16'b0000000000000000;
		15'h1046: char_row_bitmap <= 16'b0011111111000000;
		15'h1047: char_row_bitmap <= 16'b0011111111100000;
		15'h1048: char_row_bitmap <= 16'b0011000001110000;
		15'h1049: char_row_bitmap <= 16'b0011000001110000;
		15'h104a: char_row_bitmap <= 16'b0011111111100000;
		15'h104b: char_row_bitmap <= 16'b0011111111000000;
		15'h104c: char_row_bitmap <= 16'b0011000000000000;
		15'h104d: char_row_bitmap <= 16'b0011000000000000;
		15'h104e: char_row_bitmap <= 16'b0011000000000000;
		15'h104f: char_row_bitmap <= 16'b0011000000000000;
		15'h1050: char_row_bitmap <= 16'b0000000000000000;
		15'h1051: char_row_bitmap <= 16'b0000000000000000;
		15'h1052: char_row_bitmap <= 16'b0000000000000000;
		15'h1053: char_row_bitmap <= 16'b0000000000000000;
		15'h1054: char_row_bitmap <= 16'b0000000000000000;
		15'h1055: char_row_bitmap <= 16'b0000000000000000;
		15'h1056: char_row_bitmap <= 16'b0000000000000000;
		15'h1057: char_row_bitmap <= 16'b0000000000000000;
		15'h1058: char_row_bitmap <= 16'b0000000000000000;
		15'h1059: char_row_bitmap <= 16'b0000000000000000;
		15'h105a: char_row_bitmap <= 16'b0000111111000000;
		15'h105b: char_row_bitmap <= 16'b0001111111100000;
		15'h105c: char_row_bitmap <= 16'b0011100001110000;
		15'h105d: char_row_bitmap <= 16'b0011000000110000;
		15'h105e: char_row_bitmap <= 16'b0011001100110000;
		15'h105f: char_row_bitmap <= 16'b0011001110110000;
		15'h1060: char_row_bitmap <= 16'b0011000111000000;
		15'h1061: char_row_bitmap <= 16'b0011100011100000;
		15'h1062: char_row_bitmap <= 16'b0001111101110000;
		15'h1063: char_row_bitmap <= 16'b0000111100110000;
		15'h1064: char_row_bitmap <= 16'b0000000000000000;
		15'h1065: char_row_bitmap <= 16'b0000000000000000;
		15'h1066: char_row_bitmap <= 16'b0000000000000000;
		15'h1067: char_row_bitmap <= 16'b0000000000000000;
		15'h1068: char_row_bitmap <= 16'b0000000000000000;
		15'h1069: char_row_bitmap <= 16'b0000000000000000;
		15'h106a: char_row_bitmap <= 16'b0000000000000000;
		15'h106b: char_row_bitmap <= 16'b0000000000000000;
		15'h106c: char_row_bitmap <= 16'b0000000000000000;
		15'h106d: char_row_bitmap <= 16'b0000000000000000;
		15'h106e: char_row_bitmap <= 16'b0011111111000000;
		15'h106f: char_row_bitmap <= 16'b0011111111100000;
		15'h1070: char_row_bitmap <= 16'b0011000001110000;
		15'h1071: char_row_bitmap <= 16'b0011000001110000;
		15'h1072: char_row_bitmap <= 16'b0011111111100000;
		15'h1073: char_row_bitmap <= 16'b0011111111000000;
		15'h1074: char_row_bitmap <= 16'b0011011100000000;
		15'h1075: char_row_bitmap <= 16'b0011001110000000;
		15'h1076: char_row_bitmap <= 16'b0011000111000000;
		15'h1077: char_row_bitmap <= 16'b0011000011000000;
		15'h1078: char_row_bitmap <= 16'b0000000000000000;
		15'h1079: char_row_bitmap <= 16'b0000000000000000;
		15'h107a: char_row_bitmap <= 16'b0000000000000000;
		15'h107b: char_row_bitmap <= 16'b0000000000000000;
		15'h107c: char_row_bitmap <= 16'b0000000000000000;
		15'h107d: char_row_bitmap <= 16'b0000000000000000;
		15'h107e: char_row_bitmap <= 16'b0000000000000000;
		15'h107f: char_row_bitmap <= 16'b0000000000000000;
		15'h1080: char_row_bitmap <= 16'b0000000000000000;
		15'h1081: char_row_bitmap <= 16'b0000000000000000;
		15'h1082: char_row_bitmap <= 16'b0000111111110000;
		15'h1083: char_row_bitmap <= 16'b0001111111110000;
		15'h1084: char_row_bitmap <= 16'b0011100000000000;
		15'h1085: char_row_bitmap <= 16'b0011000000000000;
		15'h1086: char_row_bitmap <= 16'b0011111111110000;
		15'h1087: char_row_bitmap <= 16'b0011111111110000;
		15'h1088: char_row_bitmap <= 16'b0000000000110000;
		15'h1089: char_row_bitmap <= 16'b0000000001110000;
		15'h108a: char_row_bitmap <= 16'b0011111111100000;
		15'h108b: char_row_bitmap <= 16'b0011111111000000;
		15'h108c: char_row_bitmap <= 16'b0000000000000000;
		15'h108d: char_row_bitmap <= 16'b0000000000000000;
		15'h108e: char_row_bitmap <= 16'b0000000000000000;
		15'h108f: char_row_bitmap <= 16'b0000000000000000;
		15'h1090: char_row_bitmap <= 16'b0000000000000000;
		15'h1091: char_row_bitmap <= 16'b0000000000000000;
		15'h1092: char_row_bitmap <= 16'b0000000000000000;
		15'h1093: char_row_bitmap <= 16'b0000000000000000;
		15'h1094: char_row_bitmap <= 16'b0000000000000000;
		15'h1095: char_row_bitmap <= 16'b0000000000000000;
		15'h1096: char_row_bitmap <= 16'b0011111111110000;
		15'h1097: char_row_bitmap <= 16'b0011111111110000;
		15'h1098: char_row_bitmap <= 16'b0000001100000000;
		15'h1099: char_row_bitmap <= 16'b0000001100000000;
		15'h109a: char_row_bitmap <= 16'b0000001100000000;
		15'h109b: char_row_bitmap <= 16'b0000001100000000;
		15'h109c: char_row_bitmap <= 16'b0000001100000000;
		15'h109d: char_row_bitmap <= 16'b0000001100000000;
		15'h109e: char_row_bitmap <= 16'b0000001100000000;
		15'h109f: char_row_bitmap <= 16'b0000001100000000;
		15'h10a0: char_row_bitmap <= 16'b0000000000000000;
		15'h10a1: char_row_bitmap <= 16'b0000000000000000;
		15'h10a2: char_row_bitmap <= 16'b0000000000000000;
		15'h10a3: char_row_bitmap <= 16'b0000000000000000;
		15'h10a4: char_row_bitmap <= 16'b0000000000000000;
		15'h10a5: char_row_bitmap <= 16'b0000000000000000;
		15'h10a6: char_row_bitmap <= 16'b0000000000000000;
		15'h10a7: char_row_bitmap <= 16'b0000000000000000;
		15'h10a8: char_row_bitmap <= 16'b0000000000000000;
		15'h10a9: char_row_bitmap <= 16'b0000000000000000;
		15'h10aa: char_row_bitmap <= 16'b0011000000110000;
		15'h10ab: char_row_bitmap <= 16'b0011000000110000;
		15'h10ac: char_row_bitmap <= 16'b0011000000110000;
		15'h10ad: char_row_bitmap <= 16'b0011000000110000;
		15'h10ae: char_row_bitmap <= 16'b0011000000110000;
		15'h10af: char_row_bitmap <= 16'b0011000000110000;
		15'h10b0: char_row_bitmap <= 16'b0011000000110000;
		15'h10b1: char_row_bitmap <= 16'b0011100001110000;
		15'h10b2: char_row_bitmap <= 16'b0001111111100000;
		15'h10b3: char_row_bitmap <= 16'b0000111111000000;
		15'h10b4: char_row_bitmap <= 16'b0000000000000000;
		15'h10b5: char_row_bitmap <= 16'b0000000000000000;
		15'h10b6: char_row_bitmap <= 16'b0000000000000000;
		15'h10b7: char_row_bitmap <= 16'b0000000000000000;
		15'h10b8: char_row_bitmap <= 16'b0000000000000000;
		15'h10b9: char_row_bitmap <= 16'b0000000000000000;
		15'h10ba: char_row_bitmap <= 16'b0000000000000000;
		15'h10bb: char_row_bitmap <= 16'b0000000000000000;
		15'h10bc: char_row_bitmap <= 16'b0000000000000000;
		15'h10bd: char_row_bitmap <= 16'b0000000000000000;
		15'h10be: char_row_bitmap <= 16'b0011000000110000;
		15'h10bf: char_row_bitmap <= 16'b0011000000110000;
		15'h10c0: char_row_bitmap <= 16'b0011000000110000;
		15'h10c1: char_row_bitmap <= 16'b0011000000110000;
		15'h10c2: char_row_bitmap <= 16'b0011000000110000;
		15'h10c3: char_row_bitmap <= 16'b0011100001110000;
		15'h10c4: char_row_bitmap <= 16'b0001110011100000;
		15'h10c5: char_row_bitmap <= 16'b0000111111000000;
		15'h10c6: char_row_bitmap <= 16'b0000011110000000;
		15'h10c7: char_row_bitmap <= 16'b0000001100000000;
		15'h10c8: char_row_bitmap <= 16'b0000000000000000;
		15'h10c9: char_row_bitmap <= 16'b0000000000000000;
		15'h10ca: char_row_bitmap <= 16'b0000000000000000;
		15'h10cb: char_row_bitmap <= 16'b0000000000000000;
		15'h10cc: char_row_bitmap <= 16'b0000000000000000;
		15'h10cd: char_row_bitmap <= 16'b0000000000000000;
		15'h10ce: char_row_bitmap <= 16'b0000000000000000;
		15'h10cf: char_row_bitmap <= 16'b0000000000000000;
		15'h10d0: char_row_bitmap <= 16'b0000000000000000;
		15'h10d1: char_row_bitmap <= 16'b0000000000000000;
		15'h10d2: char_row_bitmap <= 16'b0011000000110000;
		15'h10d3: char_row_bitmap <= 16'b0011000000110000;
		15'h10d4: char_row_bitmap <= 16'b0011000000110000;
		15'h10d5: char_row_bitmap <= 16'b0011000000110000;
		15'h10d6: char_row_bitmap <= 16'b0011001100110000;
		15'h10d7: char_row_bitmap <= 16'b0011001100110000;
		15'h10d8: char_row_bitmap <= 16'b0011001100110000;
		15'h10d9: char_row_bitmap <= 16'b0011001101110000;
		15'h10da: char_row_bitmap <= 16'b0011111111100000;
		15'h10db: char_row_bitmap <= 16'b0011111111000000;
		15'h10dc: char_row_bitmap <= 16'b0000000000000000;
		15'h10dd: char_row_bitmap <= 16'b0000000000000000;
		15'h10de: char_row_bitmap <= 16'b0000000000000000;
		15'h10df: char_row_bitmap <= 16'b0000000000000000;
		15'h10e0: char_row_bitmap <= 16'b0000000000000000;
		15'h10e1: char_row_bitmap <= 16'b0000000000000000;
		15'h10e2: char_row_bitmap <= 16'b0000000000000000;
		15'h10e3: char_row_bitmap <= 16'b0000000000000000;
		15'h10e4: char_row_bitmap <= 16'b0000000000000000;
		15'h10e5: char_row_bitmap <= 16'b0000000000000000;
		15'h10e6: char_row_bitmap <= 16'b0011000000110000;
		15'h10e7: char_row_bitmap <= 16'b0011100001110000;
		15'h10e8: char_row_bitmap <= 16'b0001110011100000;
		15'h10e9: char_row_bitmap <= 16'b0000111111000000;
		15'h10ea: char_row_bitmap <= 16'b0000011110000000;
		15'h10eb: char_row_bitmap <= 16'b0000011110000000;
		15'h10ec: char_row_bitmap <= 16'b0000111111000000;
		15'h10ed: char_row_bitmap <= 16'b0001110011100000;
		15'h10ee: char_row_bitmap <= 16'b0011100001110000;
		15'h10ef: char_row_bitmap <= 16'b0011000000110000;
		15'h10f0: char_row_bitmap <= 16'b0000000000000000;
		15'h10f1: char_row_bitmap <= 16'b0000000000000000;
		15'h10f2: char_row_bitmap <= 16'b0000000000000000;
		15'h10f3: char_row_bitmap <= 16'b0000000000000000;
		15'h10f4: char_row_bitmap <= 16'b0000000000000000;
		15'h10f5: char_row_bitmap <= 16'b0000000000000000;
		15'h10f6: char_row_bitmap <= 16'b0000000000000000;
		15'h10f7: char_row_bitmap <= 16'b0000000000000000;
		15'h10f8: char_row_bitmap <= 16'b0000000000000000;
		15'h10f9: char_row_bitmap <= 16'b0000000000000000;
		15'h10fa: char_row_bitmap <= 16'b0011000000110000;
		15'h10fb: char_row_bitmap <= 16'b0011100001110000;
		15'h10fc: char_row_bitmap <= 16'b0001110011100000;
		15'h10fd: char_row_bitmap <= 16'b0000111111000000;
		15'h10fe: char_row_bitmap <= 16'b0000011110000000;
		15'h10ff: char_row_bitmap <= 16'b0000001100000000;
		15'h1100: char_row_bitmap <= 16'b0000001100000000;
		15'h1101: char_row_bitmap <= 16'b0000001100000000;
		15'h1102: char_row_bitmap <= 16'b0000001100000000;
		15'h1103: char_row_bitmap <= 16'b0000001100000000;
		15'h1104: char_row_bitmap <= 16'b0000000000000000;
		15'h1105: char_row_bitmap <= 16'b0000000000000000;
		15'h1106: char_row_bitmap <= 16'b0000000000000000;
		15'h1107: char_row_bitmap <= 16'b0000000000000000;
		15'h1108: char_row_bitmap <= 16'b0000000000000000;
		15'h1109: char_row_bitmap <= 16'b0000000000000000;
		15'h110a: char_row_bitmap <= 16'b0000000000000000;
		15'h110b: char_row_bitmap <= 16'b0000000000000000;
		15'h110c: char_row_bitmap <= 16'b0000000000000000;
		15'h110d: char_row_bitmap <= 16'b0000000000000000;
		15'h110e: char_row_bitmap <= 16'b0011111111110000;
		15'h110f: char_row_bitmap <= 16'b0011111111110000;
		15'h1110: char_row_bitmap <= 16'b0000000011100000;
		15'h1111: char_row_bitmap <= 16'b0000000111000000;
		15'h1112: char_row_bitmap <= 16'b0000001110000000;
		15'h1113: char_row_bitmap <= 16'b0000011100000000;
		15'h1114: char_row_bitmap <= 16'b0000111000000000;
		15'h1115: char_row_bitmap <= 16'b0001110000000000;
		15'h1116: char_row_bitmap <= 16'b0011111111110000;
		15'h1117: char_row_bitmap <= 16'b0011111111110000;
		15'h1118: char_row_bitmap <= 16'b0000000000000000;
		15'h1119: char_row_bitmap <= 16'b0000000000000000;
		15'h111a: char_row_bitmap <= 16'b0000000000000000;
		15'h111b: char_row_bitmap <= 16'b0000000000000000;
		15'h111c: char_row_bitmap <= 16'b0000000000000000;
		15'h111d: char_row_bitmap <= 16'b0000000000000000;
		15'h111e: char_row_bitmap <= 16'b0011000000110000;
		15'h111f: char_row_bitmap <= 16'b0011000000110000;
		15'h1120: char_row_bitmap <= 16'b0011000000110000;
		15'h1121: char_row_bitmap <= 16'b0011100001110000;
		15'h1122: char_row_bitmap <= 16'b0001100001100000;
		15'h1123: char_row_bitmap <= 16'b0001111111100000;
		15'h1124: char_row_bitmap <= 16'b0001111111100000;
		15'h1125: char_row_bitmap <= 16'b0000110011000000;
		15'h1126: char_row_bitmap <= 16'b0000110011000000;
		15'h1127: char_row_bitmap <= 16'b0000110011000000;
		15'h1128: char_row_bitmap <= 16'b0000011110000000;
		15'h1129: char_row_bitmap <= 16'b0000011110000000;
		15'h112a: char_row_bitmap <= 16'b0000001100000000;
		15'h112b: char_row_bitmap <= 16'b0000001100000000;
		15'h112c: char_row_bitmap <= 16'b0000000000000000;
		15'h112d: char_row_bitmap <= 16'b0000000000000000;
		15'h112e: char_row_bitmap <= 16'b0000000000000000;
		15'h112f: char_row_bitmap <= 16'b0000000000000000;
		15'h1130: char_row_bitmap <= 16'b0000000000000000;
		15'h1131: char_row_bitmap <= 16'b0000000000000000;
		15'h1132: char_row_bitmap <= 16'b0011111111110000;
		15'h1133: char_row_bitmap <= 16'b0011111111110000;
		15'h1134: char_row_bitmap <= 16'b0000000000110000;
		15'h1135: char_row_bitmap <= 16'b0000000000110000;
		15'h1136: char_row_bitmap <= 16'b0000000000110000;
		15'h1137: char_row_bitmap <= 16'b0000000000110000;
		15'h1138: char_row_bitmap <= 16'b0011111111110000;
		15'h1139: char_row_bitmap <= 16'b0011111111110000;
		15'h113a: char_row_bitmap <= 16'b0000000000110000;
		15'h113b: char_row_bitmap <= 16'b0000000000110000;
		15'h113c: char_row_bitmap <= 16'b0000000000110000;
		15'h113d: char_row_bitmap <= 16'b0000000000110000;
		15'h113e: char_row_bitmap <= 16'b0011111111110000;
		15'h113f: char_row_bitmap <= 16'b0011111111110000;
		15'h1140: char_row_bitmap <= 16'b0000000000000000;
		15'h1141: char_row_bitmap <= 16'b0000000000000000;
		15'h1142: char_row_bitmap <= 16'b0000000000000000;
		15'h1143: char_row_bitmap <= 16'b0000000000000000;
		15'h1144: char_row_bitmap <= 16'b0000000000000000;
		15'h1145: char_row_bitmap <= 16'b0000000000000000;
		15'h1146: char_row_bitmap <= 16'b0000000000000000;
		15'h1147: char_row_bitmap <= 16'b0000000000000000;
		15'h1148: char_row_bitmap <= 16'b0000000000000000;
		15'h1149: char_row_bitmap <= 16'b0000000000000000;
		15'h114a: char_row_bitmap <= 16'b0000000000000000;
		15'h114b: char_row_bitmap <= 16'b0000000000000000;
		15'h114c: char_row_bitmap <= 16'b0000001100000000;
		15'h114d: char_row_bitmap <= 16'b0000001100000000;
		15'h114e: char_row_bitmap <= 16'b0000011110000000;
		15'h114f: char_row_bitmap <= 16'b0000011110000000;
		15'h1150: char_row_bitmap <= 16'b0000110011000000;
		15'h1151: char_row_bitmap <= 16'b0000110011000000;
		15'h1152: char_row_bitmap <= 16'b0001100001100000;
		15'h1153: char_row_bitmap <= 16'b0001100001100000;
		15'h1154: char_row_bitmap <= 16'b0000000000000000;
		15'h1155: char_row_bitmap <= 16'b0000000000000000;
		15'h1156: char_row_bitmap <= 16'b0000000000000000;
		15'h1157: char_row_bitmap <= 16'b0000000000000000;
		15'h1158: char_row_bitmap <= 16'b0000000000000000;
		15'h1159: char_row_bitmap <= 16'b0000000000000000;
		15'h115a: char_row_bitmap <= 16'b0000000000000000;
		15'h115b: char_row_bitmap <= 16'b0000000000000000;
		15'h115c: char_row_bitmap <= 16'b0000000000000000;
		15'h115d: char_row_bitmap <= 16'b0000000000000000;
		15'h115e: char_row_bitmap <= 16'b0000000000000000;
		15'h115f: char_row_bitmap <= 16'b0000000000000000;
		15'h1160: char_row_bitmap <= 16'b0001100001100000;
		15'h1161: char_row_bitmap <= 16'b0001100001100000;
		15'h1162: char_row_bitmap <= 16'b0000110011000000;
		15'h1163: char_row_bitmap <= 16'b0000110011000000;
		15'h1164: char_row_bitmap <= 16'b0000011110000000;
		15'h1165: char_row_bitmap <= 16'b0000011110000000;
		15'h1166: char_row_bitmap <= 16'b0000001100000000;
		15'h1167: char_row_bitmap <= 16'b0000001100000000;
		15'h1168: char_row_bitmap <= 16'b0000000000000000;
		15'h1169: char_row_bitmap <= 16'b0000000000000000;
		15'h116a: char_row_bitmap <= 16'b0000000000000000;
		15'h116b: char_row_bitmap <= 16'b0000000000000000;
		15'h116c: char_row_bitmap <= 16'b0000000000000000;
		15'h116d: char_row_bitmap <= 16'b0000000000000000;
		15'h116e: char_row_bitmap <= 16'b0000000000000000;
		15'h116f: char_row_bitmap <= 16'b0000000000000000;
		15'h1170: char_row_bitmap <= 16'b0011000000000000;
		15'h1171: char_row_bitmap <= 16'b0111100001100000;
		15'h1172: char_row_bitmap <= 16'b0111100011100000;
		15'h1173: char_row_bitmap <= 16'b0011000111000000;
		15'h1174: char_row_bitmap <= 16'b0000001110000000;
		15'h1175: char_row_bitmap <= 16'b0000011100000000;
		15'h1176: char_row_bitmap <= 16'b0000111000000000;
		15'h1177: char_row_bitmap <= 16'b0001110000000000;
		15'h1178: char_row_bitmap <= 16'b0011100000000000;
		15'h1179: char_row_bitmap <= 16'b0111001100011000;
		15'h117a: char_row_bitmap <= 16'b0110011110111100;
		15'h117b: char_row_bitmap <= 16'b0000011110111100;
		15'h117c: char_row_bitmap <= 16'b0000001100011000;
		15'h117d: char_row_bitmap <= 16'b0000000000000000;
		15'h117e: char_row_bitmap <= 16'b0000000000000000;
		15'h117f: char_row_bitmap <= 16'b0000000000000000;
		15'h1180: char_row_bitmap <= 16'b0000000000000000;
		15'h1181: char_row_bitmap <= 16'b0000000000000000;
		15'h1182: char_row_bitmap <= 16'b0000000000000000;
		15'h1183: char_row_bitmap <= 16'b0000000000000000;
		15'h1184: char_row_bitmap <= 16'b0000000000000000;
		15'h1185: char_row_bitmap <= 16'b0000100100000000;
		15'h1186: char_row_bitmap <= 16'b0000110100000000;
		15'h1187: char_row_bitmap <= 16'b0000101100000000;
		15'h1188: char_row_bitmap <= 16'b0000100100000000;
		15'h1189: char_row_bitmap <= 16'b0000100100000000;
		15'h118a: char_row_bitmap <= 16'b0000000000000000;
		15'h118b: char_row_bitmap <= 16'b0000000001000000;
		15'h118c: char_row_bitmap <= 16'b0000000001000000;
		15'h118d: char_row_bitmap <= 16'b0000000001000000;
		15'h118e: char_row_bitmap <= 16'b0000000001000000;
		15'h118f: char_row_bitmap <= 16'b0000000001111000;
		15'h1190: char_row_bitmap <= 16'b0000000000000000;
		15'h1191: char_row_bitmap <= 16'b0000000000000000;
		15'h1192: char_row_bitmap <= 16'b0000000000000000;
		15'h1193: char_row_bitmap <= 16'b0000000000000000;
		15'h1194: char_row_bitmap <= 16'b0000000000000000;
		15'h1195: char_row_bitmap <= 16'b0000000000000000;
		15'h1196: char_row_bitmap <= 16'b0000000000000000;
		15'h1197: char_row_bitmap <= 16'b0000011110110000;
		15'h1198: char_row_bitmap <= 16'b0000111111110000;
		15'h1199: char_row_bitmap <= 16'b0000110001110000;
		15'h119a: char_row_bitmap <= 16'b0000110000110000;
		15'h119b: char_row_bitmap <= 16'b0000110001110000;
		15'h119c: char_row_bitmap <= 16'b0000111111110000;
		15'h119d: char_row_bitmap <= 16'b0000011110110000;
		15'h119e: char_row_bitmap <= 16'b0000000000000000;
		15'h119f: char_row_bitmap <= 16'b0000000000000000;
		15'h11a0: char_row_bitmap <= 16'b0000000000000000;
		15'h11a1: char_row_bitmap <= 16'b0000000000000000;
		15'h11a2: char_row_bitmap <= 16'b0000000000000000;
		15'h11a3: char_row_bitmap <= 16'b0000000000000000;
		15'h11a4: char_row_bitmap <= 16'b0000000000000000;
		15'h11a5: char_row_bitmap <= 16'b0000000000000000;
		15'h11a6: char_row_bitmap <= 16'b0000000000000000;
		15'h11a7: char_row_bitmap <= 16'b0000000000000000;
		15'h11a8: char_row_bitmap <= 16'b0000000000000000;
		15'h11a9: char_row_bitmap <= 16'b0000000000000000;
		15'h11aa: char_row_bitmap <= 16'b0000110000000000;
		15'h11ab: char_row_bitmap <= 16'b0000110000000000;
		15'h11ac: char_row_bitmap <= 16'b0000111111100000;
		15'h11ad: char_row_bitmap <= 16'b0000111111110000;
		15'h11ae: char_row_bitmap <= 16'b0000110000110000;
		15'h11af: char_row_bitmap <= 16'b0000110000110000;
		15'h11b0: char_row_bitmap <= 16'b0000111111110000;
		15'h11b1: char_row_bitmap <= 16'b0000111111100000;
		15'h11b2: char_row_bitmap <= 16'b0000000000000000;
		15'h11b3: char_row_bitmap <= 16'b0000000000000000;
		15'h11b4: char_row_bitmap <= 16'b0000000000000000;
		15'h11b5: char_row_bitmap <= 16'b0000000000000000;
		15'h11b6: char_row_bitmap <= 16'b0000000000000000;
		15'h11b7: char_row_bitmap <= 16'b0000000000000000;
		15'h11b8: char_row_bitmap <= 16'b0000000000000000;
		15'h11b9: char_row_bitmap <= 16'b0000000000000000;
		15'h11ba: char_row_bitmap <= 16'b0000000000000000;
		15'h11bb: char_row_bitmap <= 16'b0000000000000000;
		15'h11bc: char_row_bitmap <= 16'b0000000000000000;
		15'h11bd: char_row_bitmap <= 16'b0000000000000000;
		15'h11be: char_row_bitmap <= 16'b0000011111100000;
		15'h11bf: char_row_bitmap <= 16'b0000111111100000;
		15'h11c0: char_row_bitmap <= 16'b0000110000000000;
		15'h11c1: char_row_bitmap <= 16'b0000110000000000;
		15'h11c2: char_row_bitmap <= 16'b0000110000000000;
		15'h11c3: char_row_bitmap <= 16'b0000110000000000;
		15'h11c4: char_row_bitmap <= 16'b0000111111100000;
		15'h11c5: char_row_bitmap <= 16'b0000011111100000;
		15'h11c6: char_row_bitmap <= 16'b0000000000000000;
		15'h11c7: char_row_bitmap <= 16'b0000000000000000;
		15'h11c8: char_row_bitmap <= 16'b0000000000000000;
		15'h11c9: char_row_bitmap <= 16'b0000000000000000;
		15'h11ca: char_row_bitmap <= 16'b0000000000000000;
		15'h11cb: char_row_bitmap <= 16'b0000000000000000;
		15'h11cc: char_row_bitmap <= 16'b0000000000000000;
		15'h11cd: char_row_bitmap <= 16'b0000000000000000;
		15'h11ce: char_row_bitmap <= 16'b0000000000000000;
		15'h11cf: char_row_bitmap <= 16'b0000000000000000;
		15'h11d0: char_row_bitmap <= 16'b0000000000000000;
		15'h11d1: char_row_bitmap <= 16'b0000000000000000;
		15'h11d2: char_row_bitmap <= 16'b0000000000110000;
		15'h11d3: char_row_bitmap <= 16'b0000000000110000;
		15'h11d4: char_row_bitmap <= 16'b0000011111110000;
		15'h11d5: char_row_bitmap <= 16'b0000111111110000;
		15'h11d6: char_row_bitmap <= 16'b0000110000110000;
		15'h11d7: char_row_bitmap <= 16'b0000110000110000;
		15'h11d8: char_row_bitmap <= 16'b0000111111110000;
		15'h11d9: char_row_bitmap <= 16'b0000011111110000;
		15'h11da: char_row_bitmap <= 16'b0000000000000000;
		15'h11db: char_row_bitmap <= 16'b0000000000000000;
		15'h11dc: char_row_bitmap <= 16'b0000000000000000;
		15'h11dd: char_row_bitmap <= 16'b0000000000000000;
		15'h11de: char_row_bitmap <= 16'b0000000000000000;
		15'h11df: char_row_bitmap <= 16'b0000000000000000;
		15'h11e0: char_row_bitmap <= 16'b0000000000000000;
		15'h11e1: char_row_bitmap <= 16'b0000000000000000;
		15'h11e2: char_row_bitmap <= 16'b0000000000000000;
		15'h11e3: char_row_bitmap <= 16'b0000000000000000;
		15'h11e4: char_row_bitmap <= 16'b0000000000000000;
		15'h11e5: char_row_bitmap <= 16'b0000000000000000;
		15'h11e6: char_row_bitmap <= 16'b0000011111100000;
		15'h11e7: char_row_bitmap <= 16'b0000111111110000;
		15'h11e8: char_row_bitmap <= 16'b0000110000110000;
		15'h11e9: char_row_bitmap <= 16'b0000111111110000;
		15'h11ea: char_row_bitmap <= 16'b0000111111100000;
		15'h11eb: char_row_bitmap <= 16'b0000110000000000;
		15'h11ec: char_row_bitmap <= 16'b0000111111100000;
		15'h11ed: char_row_bitmap <= 16'b0000011111100000;
		15'h11ee: char_row_bitmap <= 16'b0000000000000000;
		15'h11ef: char_row_bitmap <= 16'b0000000000000000;
		15'h11f0: char_row_bitmap <= 16'b0000000000000000;
		15'h11f1: char_row_bitmap <= 16'b0000000000000000;
		15'h11f2: char_row_bitmap <= 16'b0000000000000000;
		15'h11f3: char_row_bitmap <= 16'b0000000000000000;
		15'h11f4: char_row_bitmap <= 16'b0000000000000000;
		15'h11f5: char_row_bitmap <= 16'b0000000000000000;
		15'h11f6: char_row_bitmap <= 16'b0000000000000000;
		15'h11f7: char_row_bitmap <= 16'b0000000000000000;
		15'h11f8: char_row_bitmap <= 16'b0000000000000000;
		15'h11f9: char_row_bitmap <= 16'b0000000000000000;
		15'h11fa: char_row_bitmap <= 16'b0000000111100000;
		15'h11fb: char_row_bitmap <= 16'b0000001111110000;
		15'h11fc: char_row_bitmap <= 16'b0000001100110000;
		15'h11fd: char_row_bitmap <= 16'b0000001100000000;
		15'h11fe: char_row_bitmap <= 16'b0000111111000000;
		15'h11ff: char_row_bitmap <= 16'b0000001100000000;
		15'h1200: char_row_bitmap <= 16'b0000001100000000;
		15'h1201: char_row_bitmap <= 16'b0000001100000000;
		15'h1202: char_row_bitmap <= 16'b0000000000000000;
		15'h1203: char_row_bitmap <= 16'b0000000000000000;
		15'h1204: char_row_bitmap <= 16'b0000000000000000;
		15'h1205: char_row_bitmap <= 16'b0000000000000000;
		15'h1206: char_row_bitmap <= 16'b0000000000000000;
		15'h1207: char_row_bitmap <= 16'b0000000000000000;
		15'h1208: char_row_bitmap <= 16'b0000000000000000;
		15'h1209: char_row_bitmap <= 16'b0000000000000000;
		15'h120a: char_row_bitmap <= 16'b0000000000000000;
		15'h120b: char_row_bitmap <= 16'b0000000000000000;
		15'h120c: char_row_bitmap <= 16'b0000000000000000;
		15'h120d: char_row_bitmap <= 16'b0000000000000000;
		15'h120e: char_row_bitmap <= 16'b0000011111100000;
		15'h120f: char_row_bitmap <= 16'b0000111111110000;
		15'h1210: char_row_bitmap <= 16'b0000110000110000;
		15'h1211: char_row_bitmap <= 16'b0000111111110000;
		15'h1212: char_row_bitmap <= 16'b0000011111110000;
		15'h1213: char_row_bitmap <= 16'b0000000000110000;
		15'h1214: char_row_bitmap <= 16'b0000110000110000;
		15'h1215: char_row_bitmap <= 16'b0000111111110000;
		15'h1216: char_row_bitmap <= 16'b0000011111100000;
		15'h1217: char_row_bitmap <= 16'b0000000000000000;
		15'h1218: char_row_bitmap <= 16'b0000000000000000;
		15'h1219: char_row_bitmap <= 16'b0000000000000000;
		15'h121a: char_row_bitmap <= 16'b0000000000000000;
		15'h121b: char_row_bitmap <= 16'b0000000000000000;
		15'h121c: char_row_bitmap <= 16'b0000000000000000;
		15'h121d: char_row_bitmap <= 16'b0000000000000000;
		15'h121e: char_row_bitmap <= 16'b0000000000000000;
		15'h121f: char_row_bitmap <= 16'b0000000000000000;
		15'h1220: char_row_bitmap <= 16'b0000000000000000;
		15'h1221: char_row_bitmap <= 16'b0000000000000000;
		15'h1222: char_row_bitmap <= 16'b0000110000000000;
		15'h1223: char_row_bitmap <= 16'b0000110000000000;
		15'h1224: char_row_bitmap <= 16'b0000110000000000;
		15'h1225: char_row_bitmap <= 16'b0000111111100000;
		15'h1226: char_row_bitmap <= 16'b0000111111110000;
		15'h1227: char_row_bitmap <= 16'b0000110000110000;
		15'h1228: char_row_bitmap <= 16'b0000110000110000;
		15'h1229: char_row_bitmap <= 16'b0000110000110000;
		15'h122a: char_row_bitmap <= 16'b0000000000000000;
		15'h122b: char_row_bitmap <= 16'b0000000000000000;
		15'h122c: char_row_bitmap <= 16'b0000000000000000;
		15'h122d: char_row_bitmap <= 16'b0000000000000000;
		15'h122e: char_row_bitmap <= 16'b0000000000000000;
		15'h122f: char_row_bitmap <= 16'b0000000000000000;
		15'h1230: char_row_bitmap <= 16'b0000000000000000;
		15'h1231: char_row_bitmap <= 16'b0000000000000000;
		15'h1232: char_row_bitmap <= 16'b0000000000000000;
		15'h1233: char_row_bitmap <= 16'b0000000000000000;
		15'h1234: char_row_bitmap <= 16'b0000000000000000;
		15'h1235: char_row_bitmap <= 16'b0000000000000000;
		15'h1236: char_row_bitmap <= 16'b0000000110000000;
		15'h1237: char_row_bitmap <= 16'b0000000110000000;
		15'h1238: char_row_bitmap <= 16'b0000000000000000;
		15'h1239: char_row_bitmap <= 16'b0000001110000000;
		15'h123a: char_row_bitmap <= 16'b0000001110000000;
		15'h123b: char_row_bitmap <= 16'b0000000110000000;
		15'h123c: char_row_bitmap <= 16'b0000000110000000;
		15'h123d: char_row_bitmap <= 16'b0000000110000000;
		15'h123e: char_row_bitmap <= 16'b0000000000000000;
		15'h123f: char_row_bitmap <= 16'b0000000000000000;
		15'h1240: char_row_bitmap <= 16'b0000000000000000;
		15'h1241: char_row_bitmap <= 16'b0000000000000000;
		15'h1242: char_row_bitmap <= 16'b0000000000000000;
		15'h1243: char_row_bitmap <= 16'b0000000000000000;
		15'h1244: char_row_bitmap <= 16'b0000000000000000;
		15'h1245: char_row_bitmap <= 16'b0000000000000000;
		15'h1246: char_row_bitmap <= 16'b0000000000000000;
		15'h1247: char_row_bitmap <= 16'b0000000000000000;
		15'h1248: char_row_bitmap <= 16'b0000000000000000;
		15'h1249: char_row_bitmap <= 16'b0000000000000000;
		15'h124a: char_row_bitmap <= 16'b0000000001100000;
		15'h124b: char_row_bitmap <= 16'b0000000001100000;
		15'h124c: char_row_bitmap <= 16'b0000000000000000;
		15'h124d: char_row_bitmap <= 16'b0000000011100000;
		15'h124e: char_row_bitmap <= 16'b0000000011100000;
		15'h124f: char_row_bitmap <= 16'b0000000001100000;
		15'h1250: char_row_bitmap <= 16'b0000011001100000;
		15'h1251: char_row_bitmap <= 16'b0000011111100000;
		15'h1252: char_row_bitmap <= 16'b0000001111000000;
		15'h1253: char_row_bitmap <= 16'b0000000000000000;
		15'h1254: char_row_bitmap <= 16'b0000000000000000;
		15'h1255: char_row_bitmap <= 16'b0000000000000000;
		15'h1256: char_row_bitmap <= 16'b0000000000000000;
		15'h1257: char_row_bitmap <= 16'b0000000000000000;
		15'h1258: char_row_bitmap <= 16'b0000000000000000;
		15'h1259: char_row_bitmap <= 16'b0000000000000000;
		15'h125a: char_row_bitmap <= 16'b0000000000000000;
		15'h125b: char_row_bitmap <= 16'b0000000000000000;
		15'h125c: char_row_bitmap <= 16'b0000000000000000;
		15'h125d: char_row_bitmap <= 16'b0000000000000000;
		15'h125e: char_row_bitmap <= 16'b0000110000000000;
		15'h125f: char_row_bitmap <= 16'b0000110011000000;
		15'h1260: char_row_bitmap <= 16'b0000110111000000;
		15'h1261: char_row_bitmap <= 16'b0000111110000000;
		15'h1262: char_row_bitmap <= 16'b0000111111000000;
		15'h1263: char_row_bitmap <= 16'b0000110011100000;
		15'h1264: char_row_bitmap <= 16'b0000110001110000;
		15'h1265: char_row_bitmap <= 16'b0000110000110000;
		15'h1266: char_row_bitmap <= 16'b0000000000000000;
		15'h1267: char_row_bitmap <= 16'b0000000000000000;
		15'h1268: char_row_bitmap <= 16'b0000000000000000;
		15'h1269: char_row_bitmap <= 16'b0000000000000000;
		15'h126a: char_row_bitmap <= 16'b0000000000000000;
		15'h126b: char_row_bitmap <= 16'b0000000000000000;
		15'h126c: char_row_bitmap <= 16'b0000000000000000;
		15'h126d: char_row_bitmap <= 16'b0000000000000000;
		15'h126e: char_row_bitmap <= 16'b0000000000000000;
		15'h126f: char_row_bitmap <= 16'b0000000000000000;
		15'h1270: char_row_bitmap <= 16'b0000000000000000;
		15'h1271: char_row_bitmap <= 16'b0000000000000000;
		15'h1272: char_row_bitmap <= 16'b0000001100000000;
		15'h1273: char_row_bitmap <= 16'b0000001100000000;
		15'h1274: char_row_bitmap <= 16'b0000001100000000;
		15'h1275: char_row_bitmap <= 16'b0000001100000000;
		15'h1276: char_row_bitmap <= 16'b0000001100000000;
		15'h1277: char_row_bitmap <= 16'b0000001100000000;
		15'h1278: char_row_bitmap <= 16'b0000001111000000;
		15'h1279: char_row_bitmap <= 16'b0000000111000000;
		15'h127a: char_row_bitmap <= 16'b0000000000000000;
		15'h127b: char_row_bitmap <= 16'b0000000000000000;
		15'h127c: char_row_bitmap <= 16'b0000000000000000;
		15'h127d: char_row_bitmap <= 16'b0000000000000000;
		15'h127e: char_row_bitmap <= 16'b0000000000000000;
		15'h127f: char_row_bitmap <= 16'b0000000000000000;
		15'h1280: char_row_bitmap <= 16'b0000000000000000;
		15'h1281: char_row_bitmap <= 16'b0000000000000000;
		15'h1282: char_row_bitmap <= 16'b0000000000000000;
		15'h1283: char_row_bitmap <= 16'b0000000000000000;
		15'h1284: char_row_bitmap <= 16'b0000000000000000;
		15'h1285: char_row_bitmap <= 16'b0000000000000000;
		15'h1286: char_row_bitmap <= 16'b0000000000000000;
		15'h1287: char_row_bitmap <= 16'b0000000000000000;
		15'h1288: char_row_bitmap <= 16'b0001111111110000;
		15'h1289: char_row_bitmap <= 16'b0001111111111000;
		15'h128a: char_row_bitmap <= 16'b0001100110011000;
		15'h128b: char_row_bitmap <= 16'b0001100110011000;
		15'h128c: char_row_bitmap <= 16'b0001100110011000;
		15'h128d: char_row_bitmap <= 16'b0001100000011000;
		15'h128e: char_row_bitmap <= 16'b0000000000000000;
		15'h128f: char_row_bitmap <= 16'b0000000000000000;
		15'h1290: char_row_bitmap <= 16'b0000000000000000;
		15'h1291: char_row_bitmap <= 16'b0000000000000000;
		15'h1292: char_row_bitmap <= 16'b0000000000000000;
		15'h1293: char_row_bitmap <= 16'b0000000000000000;
		15'h1294: char_row_bitmap <= 16'b0000000000000000;
		15'h1295: char_row_bitmap <= 16'b0000000000000000;
		15'h1296: char_row_bitmap <= 16'b0000000000000000;
		15'h1297: char_row_bitmap <= 16'b0000000000000000;
		15'h1298: char_row_bitmap <= 16'b0000000000000000;
		15'h1299: char_row_bitmap <= 16'b0000000000000000;
		15'h129a: char_row_bitmap <= 16'b0000000000000000;
		15'h129b: char_row_bitmap <= 16'b0000000000000000;
		15'h129c: char_row_bitmap <= 16'b0000111111100000;
		15'h129d: char_row_bitmap <= 16'b0000111111110000;
		15'h129e: char_row_bitmap <= 16'b0000110000110000;
		15'h129f: char_row_bitmap <= 16'b0000110000110000;
		15'h12a0: char_row_bitmap <= 16'b0000110000110000;
		15'h12a1: char_row_bitmap <= 16'b0000110000110000;
		15'h12a2: char_row_bitmap <= 16'b0000000000000000;
		15'h12a3: char_row_bitmap <= 16'b0000000000000000;
		15'h12a4: char_row_bitmap <= 16'b0000000000000000;
		15'h12a5: char_row_bitmap <= 16'b0000000000000000;
		15'h12a6: char_row_bitmap <= 16'b0000000000000000;
		15'h12a7: char_row_bitmap <= 16'b0000000000000000;
		15'h12a8: char_row_bitmap <= 16'b0000000000000000;
		15'h12a9: char_row_bitmap <= 16'b0000000000000000;
		15'h12aa: char_row_bitmap <= 16'b0000000000000000;
		15'h12ab: char_row_bitmap <= 16'b0000000000000000;
		15'h12ac: char_row_bitmap <= 16'b0000000000000000;
		15'h12ad: char_row_bitmap <= 16'b0000000000000000;
		15'h12ae: char_row_bitmap <= 16'b0000000000000000;
		15'h12af: char_row_bitmap <= 16'b0000001111000000;
		15'h12b0: char_row_bitmap <= 16'b0000011111100000;
		15'h12b1: char_row_bitmap <= 16'b0000111001110000;
		15'h12b2: char_row_bitmap <= 16'b0000110000110000;
		15'h12b3: char_row_bitmap <= 16'b0000111001110000;
		15'h12b4: char_row_bitmap <= 16'b0000011111100000;
		15'h12b5: char_row_bitmap <= 16'b0000001111000000;
		15'h12b6: char_row_bitmap <= 16'b0000000000000000;
		15'h12b7: char_row_bitmap <= 16'b0000000000000000;
		15'h12b8: char_row_bitmap <= 16'b0000000000000000;
		15'h12b9: char_row_bitmap <= 16'b0000000000000000;
		15'h12ba: char_row_bitmap <= 16'b0000000000000000;
		15'h12bb: char_row_bitmap <= 16'b0000000000000000;
		15'h12bc: char_row_bitmap <= 16'b0000000000000000;
		15'h12bd: char_row_bitmap <= 16'b0000000000000000;
		15'h12be: char_row_bitmap <= 16'b0000000000000000;
		15'h12bf: char_row_bitmap <= 16'b0000000000000000;
		15'h12c0: char_row_bitmap <= 16'b0000000000000000;
		15'h12c1: char_row_bitmap <= 16'b0000000000000000;
		15'h12c2: char_row_bitmap <= 16'b0000000000000000;
		15'h12c3: char_row_bitmap <= 16'b0000111111100000;
		15'h12c4: char_row_bitmap <= 16'b0000111111110000;
		15'h12c5: char_row_bitmap <= 16'b0000110000110000;
		15'h12c6: char_row_bitmap <= 16'b0000110000110000;
		15'h12c7: char_row_bitmap <= 16'b0000111111110000;
		15'h12c8: char_row_bitmap <= 16'b0000111111100000;
		15'h12c9: char_row_bitmap <= 16'b0000110000000000;
		15'h12ca: char_row_bitmap <= 16'b0000110000000000;
		15'h12cb: char_row_bitmap <= 16'b0000000000000000;
		15'h12cc: char_row_bitmap <= 16'b0000000000000000;
		15'h12cd: char_row_bitmap <= 16'b0000000000000000;
		15'h12ce: char_row_bitmap <= 16'b0000000000000000;
		15'h12cf: char_row_bitmap <= 16'b0000000000000000;
		15'h12d0: char_row_bitmap <= 16'b0000000000000000;
		15'h12d1: char_row_bitmap <= 16'b0000000000000000;
		15'h12d2: char_row_bitmap <= 16'b0000000000000000;
		15'h12d3: char_row_bitmap <= 16'b0000000000000000;
		15'h12d4: char_row_bitmap <= 16'b0000000000000000;
		15'h12d5: char_row_bitmap <= 16'b0000000000000000;
		15'h12d6: char_row_bitmap <= 16'b0000000000000000;
		15'h12d7: char_row_bitmap <= 16'b0000011111110000;
		15'h12d8: char_row_bitmap <= 16'b0000111111110000;
		15'h12d9: char_row_bitmap <= 16'b0000110000110000;
		15'h12da: char_row_bitmap <= 16'b0000110000110000;
		15'h12db: char_row_bitmap <= 16'b0000111111110000;
		15'h12dc: char_row_bitmap <= 16'b0000011111110000;
		15'h12dd: char_row_bitmap <= 16'b0000000000110000;
		15'h12de: char_row_bitmap <= 16'b0000000000110000;
		15'h12df: char_row_bitmap <= 16'b0000000000000000;
		15'h12e0: char_row_bitmap <= 16'b0000000000000000;
		15'h12e1: char_row_bitmap <= 16'b0000000000000000;
		15'h12e2: char_row_bitmap <= 16'b0000000000000000;
		15'h12e3: char_row_bitmap <= 16'b0000000000000000;
		15'h12e4: char_row_bitmap <= 16'b0000000000000000;
		15'h12e5: char_row_bitmap <= 16'b0000000000000000;
		15'h12e6: char_row_bitmap <= 16'b0000000000000000;
		15'h12e7: char_row_bitmap <= 16'b0000000000000000;
		15'h12e8: char_row_bitmap <= 16'b0000000000000000;
		15'h12e9: char_row_bitmap <= 16'b0000000000000000;
		15'h12ea: char_row_bitmap <= 16'b0000000000000000;
		15'h12eb: char_row_bitmap <= 16'b0000110111000000;
		15'h12ec: char_row_bitmap <= 16'b0000111111100000;
		15'h12ed: char_row_bitmap <= 16'b0000111001100000;
		15'h12ee: char_row_bitmap <= 16'b0000110000000000;
		15'h12ef: char_row_bitmap <= 16'b0000110000000000;
		15'h12f0: char_row_bitmap <= 16'b0000110000000000;
		15'h12f1: char_row_bitmap <= 16'b0000110000000000;
		15'h12f2: char_row_bitmap <= 16'b0000000000000000;
		15'h12f3: char_row_bitmap <= 16'b0000000000000000;
		15'h12f4: char_row_bitmap <= 16'b0000000000000000;
		15'h12f5: char_row_bitmap <= 16'b0000000000000000;
		15'h12f6: char_row_bitmap <= 16'b0000000000000000;
		15'h12f7: char_row_bitmap <= 16'b0000000000000000;
		15'h12f8: char_row_bitmap <= 16'b0000000000000000;
		15'h12f9: char_row_bitmap <= 16'b0000000000000000;
		15'h12fa: char_row_bitmap <= 16'b0000000000000000;
		15'h12fb: char_row_bitmap <= 16'b0000000000000000;
		15'h12fc: char_row_bitmap <= 16'b0000000000000000;
		15'h12fd: char_row_bitmap <= 16'b0000000000000000;
		15'h12fe: char_row_bitmap <= 16'b0000011111000000;
		15'h12ff: char_row_bitmap <= 16'b0000111111100000;
		15'h1300: char_row_bitmap <= 16'b0000110000000000;
		15'h1301: char_row_bitmap <= 16'b0000111111000000;
		15'h1302: char_row_bitmap <= 16'b0000011111100000;
		15'h1303: char_row_bitmap <= 16'b0000000001100000;
		15'h1304: char_row_bitmap <= 16'b0000111111100000;
		15'h1305: char_row_bitmap <= 16'b0000011111000000;
		15'h1306: char_row_bitmap <= 16'b0000000000000000;
		15'h1307: char_row_bitmap <= 16'b0000000000000000;
		15'h1308: char_row_bitmap <= 16'b0000000000000000;
		15'h1309: char_row_bitmap <= 16'b0000000000000000;
		15'h130a: char_row_bitmap <= 16'b0000000000000000;
		15'h130b: char_row_bitmap <= 16'b0000000000000000;
		15'h130c: char_row_bitmap <= 16'b0000000000000000;
		15'h130d: char_row_bitmap <= 16'b0000000000000000;
		15'h130e: char_row_bitmap <= 16'b0000000000000000;
		15'h130f: char_row_bitmap <= 16'b0000000000000000;
		15'h1310: char_row_bitmap <= 16'b0000000000000000;
		15'h1311: char_row_bitmap <= 16'b0000000000000000;
		15'h1312: char_row_bitmap <= 16'b0000001100000000;
		15'h1313: char_row_bitmap <= 16'b0000001100000000;
		15'h1314: char_row_bitmap <= 16'b0000111111000000;
		15'h1315: char_row_bitmap <= 16'b0000111111000000;
		15'h1316: char_row_bitmap <= 16'b0000001100000000;
		15'h1317: char_row_bitmap <= 16'b0000001100000000;
		15'h1318: char_row_bitmap <= 16'b0000001111000000;
		15'h1319: char_row_bitmap <= 16'b0000000111000000;
		15'h131a: char_row_bitmap <= 16'b0000000000000000;
		15'h131b: char_row_bitmap <= 16'b0000000000000000;
		15'h131c: char_row_bitmap <= 16'b0000000000000000;
		15'h131d: char_row_bitmap <= 16'b0000000000000000;
		15'h131e: char_row_bitmap <= 16'b0000000000000000;
		15'h131f: char_row_bitmap <= 16'b0000000000000000;
		15'h1320: char_row_bitmap <= 16'b0000000000000000;
		15'h1321: char_row_bitmap <= 16'b0000000000000000;
		15'h1322: char_row_bitmap <= 16'b0000000000000000;
		15'h1323: char_row_bitmap <= 16'b0000000000000000;
		15'h1324: char_row_bitmap <= 16'b0000000000000000;
		15'h1325: char_row_bitmap <= 16'b0000000000000000;
		15'h1326: char_row_bitmap <= 16'b0000000000000000;
		15'h1327: char_row_bitmap <= 16'b0000110000110000;
		15'h1328: char_row_bitmap <= 16'b0000110000110000;
		15'h1329: char_row_bitmap <= 16'b0000110000110000;
		15'h132a: char_row_bitmap <= 16'b0000110000110000;
		15'h132b: char_row_bitmap <= 16'b0000110000110000;
		15'h132c: char_row_bitmap <= 16'b0000111111110000;
		15'h132d: char_row_bitmap <= 16'b0000011111100000;
		15'h132e: char_row_bitmap <= 16'b0000000000000000;
		15'h132f: char_row_bitmap <= 16'b0000000000000000;
		15'h1330: char_row_bitmap <= 16'b0000000000000000;
		15'h1331: char_row_bitmap <= 16'b0000000000000000;
		15'h1332: char_row_bitmap <= 16'b0000000000000000;
		15'h1333: char_row_bitmap <= 16'b0000000000000000;
		15'h1334: char_row_bitmap <= 16'b0000000000000000;
		15'h1335: char_row_bitmap <= 16'b0000000000000000;
		15'h1336: char_row_bitmap <= 16'b0000000000000000;
		15'h1337: char_row_bitmap <= 16'b0000000000000000;
		15'h1338: char_row_bitmap <= 16'b0000000000000000;
		15'h1339: char_row_bitmap <= 16'b0000000000000000;
		15'h133a: char_row_bitmap <= 16'b0000000000000000;
		15'h133b: char_row_bitmap <= 16'b0000110000110000;
		15'h133c: char_row_bitmap <= 16'b0000110000110000;
		15'h133d: char_row_bitmap <= 16'b0000110000110000;
		15'h133e: char_row_bitmap <= 16'b0000111001110000;
		15'h133f: char_row_bitmap <= 16'b0000011111100000;
		15'h1340: char_row_bitmap <= 16'b0000001111000000;
		15'h1341: char_row_bitmap <= 16'b0000000110000000;
		15'h1342: char_row_bitmap <= 16'b0000000000000000;
		15'h1343: char_row_bitmap <= 16'b0000000000000000;
		15'h1344: char_row_bitmap <= 16'b0000000000000000;
		15'h1345: char_row_bitmap <= 16'b0000000000000000;
		15'h1346: char_row_bitmap <= 16'b0000000000000000;
		15'h1347: char_row_bitmap <= 16'b0000000000000000;
		15'h1348: char_row_bitmap <= 16'b0000000000000000;
		15'h1349: char_row_bitmap <= 16'b0000000000000000;
		15'h134a: char_row_bitmap <= 16'b0000000000000000;
		15'h134b: char_row_bitmap <= 16'b0000000000000000;
		15'h134c: char_row_bitmap <= 16'b0000000000000000;
		15'h134d: char_row_bitmap <= 16'b0000000000000000;
		15'h134e: char_row_bitmap <= 16'b0000000000000000;
		15'h134f: char_row_bitmap <= 16'b0001100000011000;
		15'h1350: char_row_bitmap <= 16'b0001100000011000;
		15'h1351: char_row_bitmap <= 16'b0001100110011000;
		15'h1352: char_row_bitmap <= 16'b0001100110011000;
		15'h1353: char_row_bitmap <= 16'b0001110110111000;
		15'h1354: char_row_bitmap <= 16'b0000111111110000;
		15'h1355: char_row_bitmap <= 16'b0000011001100000;
		15'h1356: char_row_bitmap <= 16'b0000000000000000;
		15'h1357: char_row_bitmap <= 16'b0000000000000000;
		15'h1358: char_row_bitmap <= 16'b0000000000000000;
		15'h1359: char_row_bitmap <= 16'b0000000000000000;
		15'h135a: char_row_bitmap <= 16'b0000000000000000;
		15'h135b: char_row_bitmap <= 16'b0000000000000000;
		15'h135c: char_row_bitmap <= 16'b0000000000000000;
		15'h135d: char_row_bitmap <= 16'b0000000000000000;
		15'h135e: char_row_bitmap <= 16'b0000000000000000;
		15'h135f: char_row_bitmap <= 16'b0000000000000000;
		15'h1360: char_row_bitmap <= 16'b0000000000000000;
		15'h1361: char_row_bitmap <= 16'b0000000000000000;
		15'h1362: char_row_bitmap <= 16'b0000000000000000;
		15'h1363: char_row_bitmap <= 16'b0000110000110000;
		15'h1364: char_row_bitmap <= 16'b0000111001110000;
		15'h1365: char_row_bitmap <= 16'b0000011111100000;
		15'h1366: char_row_bitmap <= 16'b0000001111000000;
		15'h1367: char_row_bitmap <= 16'b0000011111100000;
		15'h1368: char_row_bitmap <= 16'b0000111001110000;
		15'h1369: char_row_bitmap <= 16'b0000110000110000;
		15'h136a: char_row_bitmap <= 16'b0000000000000000;
		15'h136b: char_row_bitmap <= 16'b0000000000000000;
		15'h136c: char_row_bitmap <= 16'b0000000000000000;
		15'h136d: char_row_bitmap <= 16'b0000000000000000;
		15'h136e: char_row_bitmap <= 16'b0000000000000000;
		15'h136f: char_row_bitmap <= 16'b0000000000000000;
		15'h1370: char_row_bitmap <= 16'b0000000000000000;
		15'h1371: char_row_bitmap <= 16'b0000000000000000;
		15'h1372: char_row_bitmap <= 16'b0000000000000000;
		15'h1373: char_row_bitmap <= 16'b0000000000000000;
		15'h1374: char_row_bitmap <= 16'b0000000000000000;
		15'h1375: char_row_bitmap <= 16'b0000000000000000;
		15'h1376: char_row_bitmap <= 16'b0000011001100000;
		15'h1377: char_row_bitmap <= 16'b0000011001100000;
		15'h1378: char_row_bitmap <= 16'b0000011101100000;
		15'h1379: char_row_bitmap <= 16'b0000001111100000;
		15'h137a: char_row_bitmap <= 16'b0000000111100000;
		15'h137b: char_row_bitmap <= 16'b0000000001100000;
		15'h137c: char_row_bitmap <= 16'b0000011001100000;
		15'h137d: char_row_bitmap <= 16'b0000011111100000;
		15'h137e: char_row_bitmap <= 16'b0000001111000000;
		15'h137f: char_row_bitmap <= 16'b0000000000000000;
		15'h1380: char_row_bitmap <= 16'b0000000000000000;
		15'h1381: char_row_bitmap <= 16'b0000000000000000;
		15'h1382: char_row_bitmap <= 16'b0000000000000000;
		15'h1383: char_row_bitmap <= 16'b0000000000000000;
		15'h1384: char_row_bitmap <= 16'b0000000000000000;
		15'h1385: char_row_bitmap <= 16'b0000000000000000;
		15'h1386: char_row_bitmap <= 16'b0000000000000000;
		15'h1387: char_row_bitmap <= 16'b0000000000000000;
		15'h1388: char_row_bitmap <= 16'b0000000000000000;
		15'h1389: char_row_bitmap <= 16'b0000000000000000;
		15'h138a: char_row_bitmap <= 16'b0000111111100000;
		15'h138b: char_row_bitmap <= 16'b0000111111100000;
		15'h138c: char_row_bitmap <= 16'b0000000011100000;
		15'h138d: char_row_bitmap <= 16'b0000000111000000;
		15'h138e: char_row_bitmap <= 16'b0000001110000000;
		15'h138f: char_row_bitmap <= 16'b0000011100000000;
		15'h1390: char_row_bitmap <= 16'b0000111111100000;
		15'h1391: char_row_bitmap <= 16'b0000111111100000;
		15'h1392: char_row_bitmap <= 16'b0000000000000000;
		15'h1393: char_row_bitmap <= 16'b0000000000000000;
		15'h1394: char_row_bitmap <= 16'b0000000000000000;
		15'h1395: char_row_bitmap <= 16'b0000000000000000;
		15'h1396: char_row_bitmap <= 16'b0000000000000000;
		15'h1397: char_row_bitmap <= 16'b0000000000000000;
		15'h1398: char_row_bitmap <= 16'b0000000000000000;
		15'h1399: char_row_bitmap <= 16'b0000000000000000;
		15'h139a: char_row_bitmap <= 16'b0000000000000000;
		15'h139b: char_row_bitmap <= 16'b0000000000000000;
		15'h139c: char_row_bitmap <= 16'b0000000000000000;
		15'h139d: char_row_bitmap <= 16'b0000000000000000;
		15'h139e: char_row_bitmap <= 16'b0000000000000000;
		15'h139f: char_row_bitmap <= 16'b0000000000000000;
		15'h13a0: char_row_bitmap <= 16'b0000000000000000;
		15'h13a1: char_row_bitmap <= 16'b0000000000000000;
		15'h13a2: char_row_bitmap <= 16'b0000000000000000;
		15'h13a3: char_row_bitmap <= 16'b0000000000000000;
		15'h13a4: char_row_bitmap <= 16'b0000000000000000;
		15'h13a5: char_row_bitmap <= 16'b0000000000000000;
		15'h13a6: char_row_bitmap <= 16'b0000000000000000;
		15'h13a7: char_row_bitmap <= 16'b0000000000000000;
		15'h13a8: char_row_bitmap <= 16'b0000000000000000;
		15'h13a9: char_row_bitmap <= 16'b0000000000000000;
		15'h13aa: char_row_bitmap <= 16'b0000000000000000;
		15'h13ab: char_row_bitmap <= 16'b0000000000000000;
		15'h13ac: char_row_bitmap <= 16'b0000000000000000;
		15'h13ad: char_row_bitmap <= 16'b0000000000000000;
		15'h13ae: char_row_bitmap <= 16'b0000000000000000;
		15'h13af: char_row_bitmap <= 16'b0000000000000000;
		15'h13b0: char_row_bitmap <= 16'b0000000000000000;
		15'h13b1: char_row_bitmap <= 16'b0000000000000000;
		15'h13b2: char_row_bitmap <= 16'b0000000000000000;
		15'h13b3: char_row_bitmap <= 16'b0000000000000000;
		15'h13b4: char_row_bitmap <= 16'b0000000000000000;
		15'h13b5: char_row_bitmap <= 16'b0000000000000000;
		15'h13b6: char_row_bitmap <= 16'b0000000000000000;
		15'h13b7: char_row_bitmap <= 16'b0000000000000000;
		15'h13b8: char_row_bitmap <= 16'b0000000000000000;
		15'h13b9: char_row_bitmap <= 16'b0000000000000000;
		15'h13ba: char_row_bitmap <= 16'b0000000000000000;
		15'h13bb: char_row_bitmap <= 16'b0000000000000000;
		15'h13bc: char_row_bitmap <= 16'b0000000000000000;
		15'h13bd: char_row_bitmap <= 16'b0000000000000000;
		15'h13be: char_row_bitmap <= 16'b0000000000000000;
		15'h13bf: char_row_bitmap <= 16'b0000000000000000;
		15'h13c0: char_row_bitmap <= 16'b0000000000000000;
		15'h13c1: char_row_bitmap <= 16'b0000000000000000;
		15'h13c2: char_row_bitmap <= 16'b0000000000000000;
		15'h13c3: char_row_bitmap <= 16'b0000000000000000;
		15'h13c4: char_row_bitmap <= 16'b0000000000000000;
		15'h13c5: char_row_bitmap <= 16'b0000000000000000;
		15'h13c6: char_row_bitmap <= 16'b0000000000000000;
		15'h13c7: char_row_bitmap <= 16'b0000000000000000;
		15'h13c8: char_row_bitmap <= 16'b0000000000000000;
		15'h13c9: char_row_bitmap <= 16'b0000000000000000;
		15'h13ca: char_row_bitmap <= 16'b0000000000000000;
		15'h13cb: char_row_bitmap <= 16'b0000000000000000;
		15'h13cc: char_row_bitmap <= 16'b0000000000000000;
		15'h13cd: char_row_bitmap <= 16'b0000000000000000;
		15'h13ce: char_row_bitmap <= 16'b0000000000000000;
		15'h13cf: char_row_bitmap <= 16'b0000000000000000;
		15'h13d0: char_row_bitmap <= 16'b0000000000000000;
		15'h13d1: char_row_bitmap <= 16'b0000000000000000;
		15'h13d2: char_row_bitmap <= 16'b0000000000000000;
		15'h13d3: char_row_bitmap <= 16'b0000000000000000;
		15'h13d4: char_row_bitmap <= 16'b0000000000000000;
		15'h13d5: char_row_bitmap <= 16'b0000000000000000;
		15'h13d6: char_row_bitmap <= 16'b0000000000000000;
		15'h13d7: char_row_bitmap <= 16'b0000000000000000;
		15'h13d8: char_row_bitmap <= 16'b0000000000000000;
		15'h13d9: char_row_bitmap <= 16'b0000000000000000;
		15'h13da: char_row_bitmap <= 16'b0000000000000000;
		15'h13db: char_row_bitmap <= 16'b0000000000000000;
		15'h13dc: char_row_bitmap <= 16'b0000000000000000;
		15'h13dd: char_row_bitmap <= 16'b0000000000000000;
		15'h13de: char_row_bitmap <= 16'b0000000000000000;
		15'h13df: char_row_bitmap <= 16'b0000000000000000;
		15'h13e0: char_row_bitmap <= 16'b0000000000000000;
		15'h13e1: char_row_bitmap <= 16'b0000000000000000;
		15'h13e2: char_row_bitmap <= 16'b0000000000000000;
		15'h13e3: char_row_bitmap <= 16'b0000000000000000;
		15'h13e4: char_row_bitmap <= 16'b0000000000000000;
		15'h13e5: char_row_bitmap <= 16'b0000000000000000;
		15'h13e6: char_row_bitmap <= 16'b0000000000000000;
		15'h13e7: char_row_bitmap <= 16'b0000000000000000;
		15'h13e8: char_row_bitmap <= 16'b0000000000000000;
		15'h13e9: char_row_bitmap <= 16'b0000000000000000;
		15'h13ea: char_row_bitmap <= 16'b0000000000000000;
		15'h13eb: char_row_bitmap <= 16'b0000000000000000;
		15'h13ec: char_row_bitmap <= 16'b0000000000000000;
		15'h13ed: char_row_bitmap <= 16'b0000000000000000;
		15'h13ee: char_row_bitmap <= 16'b0000000000000000;
		15'h13ef: char_row_bitmap <= 16'b0000000000000000;
		15'h13f0: char_row_bitmap <= 16'b0000000000000000;
		15'h13f1: char_row_bitmap <= 16'b0000000000000000;
		15'h13f2: char_row_bitmap <= 16'b0000000000000000;
		15'h13f3: char_row_bitmap <= 16'b0000000000000000;
		15'h13f4: char_row_bitmap <= 16'b0000000000000000;
		15'h13f5: char_row_bitmap <= 16'b0000000000000000;
		15'h13f6: char_row_bitmap <= 16'b0000000000000000;
		15'h13f7: char_row_bitmap <= 16'b0000000000000000;
		15'h13f8: char_row_bitmap <= 16'b0000000000000000;
		15'h13f9: char_row_bitmap <= 16'b0000000000000000;
		15'h13fa: char_row_bitmap <= 16'b0000000000000000;
		15'h13fb: char_row_bitmap <= 16'b0000000000000000;
		15'h13fc: char_row_bitmap <= 16'b0000000000000000;
		15'h13fd: char_row_bitmap <= 16'b0000000000000000;
		15'h13fe: char_row_bitmap <= 16'b0000000000000000;
		15'h13ff: char_row_bitmap <= 16'b0000000000000000;
		15'h1400: char_row_bitmap <= 16'b0000000000000000;
		15'h1401: char_row_bitmap <= 16'b0000000000000000;
		15'h1402: char_row_bitmap <= 16'b0000000000000000;
		15'h1403: char_row_bitmap <= 16'b0000000000000000;
		15'h1404: char_row_bitmap <= 16'b0000000000000000;
		15'h1405: char_row_bitmap <= 16'b0000000000000000;
		15'h1406: char_row_bitmap <= 16'b0000000000000000;
		15'h1407: char_row_bitmap <= 16'b0000000000000000;
		15'h1408: char_row_bitmap <= 16'b0000000000000000;
		15'h1409: char_row_bitmap <= 16'b0000000000000000;
		15'h140a: char_row_bitmap <= 16'b0000000000000000;
		15'h140b: char_row_bitmap <= 16'b0000000000000000;
		15'h140c: char_row_bitmap <= 16'b0000000000000000;
		15'h140d: char_row_bitmap <= 16'b0000000000000000;
		15'h140e: char_row_bitmap <= 16'b0000000000000000;
		15'h140f: char_row_bitmap <= 16'b0000000000000000;
		15'h1410: char_row_bitmap <= 16'b0000000000000000;
		15'h1411: char_row_bitmap <= 16'b0000000000000000;
		15'h1412: char_row_bitmap <= 16'b0000000000000000;
		15'h1413: char_row_bitmap <= 16'b0000000000000000;
		15'h1414: char_row_bitmap <= 16'b0000000000000000;
		15'h1415: char_row_bitmap <= 16'b0000000000000000;
		15'h1416: char_row_bitmap <= 16'b0000000000000000;
		15'h1417: char_row_bitmap <= 16'b0000000000000000;
		15'h1418: char_row_bitmap <= 16'b0000000000000000;
		15'h1419: char_row_bitmap <= 16'b0000000000000000;
		15'h141a: char_row_bitmap <= 16'b0000000000000000;
		15'h141b: char_row_bitmap <= 16'b0000000000000000;
		15'h141c: char_row_bitmap <= 16'b0000000000000000;
		15'h141d: char_row_bitmap <= 16'b0000000000000000;
		15'h141e: char_row_bitmap <= 16'b0000000000000000;
		15'h141f: char_row_bitmap <= 16'b0000000000000000;
		15'h1420: char_row_bitmap <= 16'b0000000000000000;
		15'h1421: char_row_bitmap <= 16'b0000000000000000;
		15'h1422: char_row_bitmap <= 16'b0000000000000000;
		15'h1423: char_row_bitmap <= 16'b0000000000000000;
		15'h1424: char_row_bitmap <= 16'b0000000000000000;
		15'h1425: char_row_bitmap <= 16'b0000000000000000;
		15'h1426: char_row_bitmap <= 16'b0000000000000000;
		15'h1427: char_row_bitmap <= 16'b0000000000000000;
		15'h1428: char_row_bitmap <= 16'b0000000000000000;
		15'h1429: char_row_bitmap <= 16'b0000000000000000;
		15'h142a: char_row_bitmap <= 16'b0000000000000000;
		15'h142b: char_row_bitmap <= 16'b0000000000000000;
		15'h142c: char_row_bitmap <= 16'b0000000000000000;
		15'h142d: char_row_bitmap <= 16'b0000000000000000;
		15'h142e: char_row_bitmap <= 16'b0000000000000000;
		15'h142f: char_row_bitmap <= 16'b0000000000000000;
		15'h1430: char_row_bitmap <= 16'b0000000000000000;
		15'h1431: char_row_bitmap <= 16'b0000000000000000;
		15'h1432: char_row_bitmap <= 16'b0000000000000000;
		15'h1433: char_row_bitmap <= 16'b0000000000000000;
		15'h1434: char_row_bitmap <= 16'b0000000000000000;
		15'h1435: char_row_bitmap <= 16'b0000000000000000;
		15'h1436: char_row_bitmap <= 16'b0000000000000000;
		15'h1437: char_row_bitmap <= 16'b0000000000000000;
		15'h1438: char_row_bitmap <= 16'b0000000000000000;
		15'h1439: char_row_bitmap <= 16'b0000000000000000;
		15'h143a: char_row_bitmap <= 16'b0000000000000000;
		15'h143b: char_row_bitmap <= 16'b0000000000000000;
		15'h143c: char_row_bitmap <= 16'b0000000000000000;
		15'h143d: char_row_bitmap <= 16'b0000000000000000;
		15'h143e: char_row_bitmap <= 16'b0000000000000000;
		15'h143f: char_row_bitmap <= 16'b0000000000000000;
		15'h1440: char_row_bitmap <= 16'b0000000000000000;
		15'h1441: char_row_bitmap <= 16'b0000000000000000;
		15'h1442: char_row_bitmap <= 16'b0000000000000000;
		15'h1443: char_row_bitmap <= 16'b0000000000000000;
		15'h1444: char_row_bitmap <= 16'b0000000000000000;
		15'h1445: char_row_bitmap <= 16'b0000000000000000;
		15'h1446: char_row_bitmap <= 16'b0000000000000000;
		15'h1447: char_row_bitmap <= 16'b0000000000000000;
		15'h1448: char_row_bitmap <= 16'b0000000000000000;
		15'h1449: char_row_bitmap <= 16'b0000000000000000;
		15'h144a: char_row_bitmap <= 16'b0000000000000000;
		15'h144b: char_row_bitmap <= 16'b0000000000000000;
		15'h144c: char_row_bitmap <= 16'b0000000000000000;
		15'h144d: char_row_bitmap <= 16'b0000000000000000;
		15'h144e: char_row_bitmap <= 16'b0000000000000000;
		15'h144f: char_row_bitmap <= 16'b0000000000000000;
		15'h1450: char_row_bitmap <= 16'b0000000000000000;
		15'h1451: char_row_bitmap <= 16'b0000000000000000;
		15'h1452: char_row_bitmap <= 16'b0000000000000000;
		15'h1453: char_row_bitmap <= 16'b0000000000000000;
		15'h1454: char_row_bitmap <= 16'b0000000000000000;
		15'h1455: char_row_bitmap <= 16'b0000000000000000;
		15'h1456: char_row_bitmap <= 16'b0000000000000000;
		15'h1457: char_row_bitmap <= 16'b0000000000000000;
		15'h1458: char_row_bitmap <= 16'b0000000000000000;
		15'h1459: char_row_bitmap <= 16'b0000000000000000;
		15'h145a: char_row_bitmap <= 16'b0000000000000000;
		15'h145b: char_row_bitmap <= 16'b0000000000000000;
		15'h145c: char_row_bitmap <= 16'b0000000000000000;
		15'h145d: char_row_bitmap <= 16'b0000000000000000;
		15'h145e: char_row_bitmap <= 16'b0000000000000000;
		15'h145f: char_row_bitmap <= 16'b0000000000000000;
		15'h1460: char_row_bitmap <= 16'b0000000000000000;
		15'h1461: char_row_bitmap <= 16'b0000000000000000;
		15'h1462: char_row_bitmap <= 16'b0000000000000000;
		15'h1463: char_row_bitmap <= 16'b0000000000000000;
		15'h1464: char_row_bitmap <= 16'b0000000000000000;
		15'h1465: char_row_bitmap <= 16'b0000000000000000;
		15'h1466: char_row_bitmap <= 16'b0000000000000000;
		15'h1467: char_row_bitmap <= 16'b0000000000000000;
		15'h1468: char_row_bitmap <= 16'b0000000000000000;
		15'h1469: char_row_bitmap <= 16'b0000000000000000;
		15'h146a: char_row_bitmap <= 16'b0000000000000000;
		15'h146b: char_row_bitmap <= 16'b0000000000000000;
		15'h146c: char_row_bitmap <= 16'b0000000000000000;
		15'h146d: char_row_bitmap <= 16'b0000000000000000;
		15'h146e: char_row_bitmap <= 16'b0000000000000000;
		15'h146f: char_row_bitmap <= 16'b0000000000000000;
		15'h1470: char_row_bitmap <= 16'b0000000000000000;
		15'h1471: char_row_bitmap <= 16'b0000000000000000;
		15'h1472: char_row_bitmap <= 16'b0000000000000000;
		15'h1473: char_row_bitmap <= 16'b0000000000000000;
		15'h1474: char_row_bitmap <= 16'b0000000000000000;
		15'h1475: char_row_bitmap <= 16'b0000000000000000;
		15'h1476: char_row_bitmap <= 16'b0000000000000000;
		15'h1477: char_row_bitmap <= 16'b0000000000000000;
		15'h1478: char_row_bitmap <= 16'b0000000000000000;
		15'h1479: char_row_bitmap <= 16'b0000000000000000;
		15'h147a: char_row_bitmap <= 16'b0000000000000000;
		15'h147b: char_row_bitmap <= 16'b0000000000000000;
		15'h147c: char_row_bitmap <= 16'b0000000000000000;
		15'h147d: char_row_bitmap <= 16'b0000000000000000;
		15'h147e: char_row_bitmap <= 16'b0000000000000000;
		15'h147f: char_row_bitmap <= 16'b0000000000000000;
		15'h1480: char_row_bitmap <= 16'b0000000000000000;
		15'h1481: char_row_bitmap <= 16'b0000000000000000;
		15'h1482: char_row_bitmap <= 16'b0000000000000000;
		15'h1483: char_row_bitmap <= 16'b0000000000000000;
		15'h1484: char_row_bitmap <= 16'b0000000000000000;
		15'h1485: char_row_bitmap <= 16'b0000000000000000;
		15'h1486: char_row_bitmap <= 16'b0000000000000000;
		15'h1487: char_row_bitmap <= 16'b0000000000000000;
		15'h1488: char_row_bitmap <= 16'b0000000000000000;
		15'h1489: char_row_bitmap <= 16'b0000000000000000;
		15'h148a: char_row_bitmap <= 16'b0000000000000000;
		15'h148b: char_row_bitmap <= 16'b0000000000000000;
		15'h148c: char_row_bitmap <= 16'b0000000000000000;
		15'h148d: char_row_bitmap <= 16'b0000000000000000;
		15'h148e: char_row_bitmap <= 16'b0000000000000000;
		15'h148f: char_row_bitmap <= 16'b0000000000000000;
		15'h1490: char_row_bitmap <= 16'b0000000000000000;
		15'h1491: char_row_bitmap <= 16'b0000000000000000;
		15'h1492: char_row_bitmap <= 16'b0000000000000000;
		15'h1493: char_row_bitmap <= 16'b0000000000000000;
		15'h1494: char_row_bitmap <= 16'b0000000000000000;
		15'h1495: char_row_bitmap <= 16'b0000000000000000;
		15'h1496: char_row_bitmap <= 16'b0000000000000000;
		15'h1497: char_row_bitmap <= 16'b0000000000000000;
		15'h1498: char_row_bitmap <= 16'b0000000000000000;
		15'h1499: char_row_bitmap <= 16'b0000000000000000;
		15'h149a: char_row_bitmap <= 16'b0000000000000000;
		15'h149b: char_row_bitmap <= 16'b0000000000000000;
		15'h149c: char_row_bitmap <= 16'b0000000000000000;
		15'h149d: char_row_bitmap <= 16'b0000000000000000;
		15'h149e: char_row_bitmap <= 16'b0000000000000000;
		15'h149f: char_row_bitmap <= 16'b0000000000000000;
		15'h14a0: char_row_bitmap <= 16'b0000000000000000;
		15'h14a1: char_row_bitmap <= 16'b0000000000000000;
		15'h14a2: char_row_bitmap <= 16'b0000000000000000;
		15'h14a3: char_row_bitmap <= 16'b0000000000000000;
		15'h14a4: char_row_bitmap <= 16'b0000000000000000;
		15'h14a5: char_row_bitmap <= 16'b0000000000000000;
		15'h14a6: char_row_bitmap <= 16'b0000000000000000;
		15'h14a7: char_row_bitmap <= 16'b0000000000000000;
		15'h14a8: char_row_bitmap <= 16'b0000000000000000;
		15'h14a9: char_row_bitmap <= 16'b0000000000000000;
		15'h14aa: char_row_bitmap <= 16'b0000000000000000;
		15'h14ab: char_row_bitmap <= 16'b0000000000000000;
		15'h14ac: char_row_bitmap <= 16'b0000000000000000;
		15'h14ad: char_row_bitmap <= 16'b0000000000000000;
		15'h14ae: char_row_bitmap <= 16'b0000000000000000;
		15'h14af: char_row_bitmap <= 16'b0000000000000000;
		15'h14b0: char_row_bitmap <= 16'b0000000000000000;
		15'h14b1: char_row_bitmap <= 16'b0000000000000000;
		15'h14b2: char_row_bitmap <= 16'b0000000000000000;
		15'h14b3: char_row_bitmap <= 16'b0000000000000000;
		15'h14b4: char_row_bitmap <= 16'b0000000000000000;
		15'h14b5: char_row_bitmap <= 16'b0000000000000000;
		15'h14b6: char_row_bitmap <= 16'b0000000000000000;
		15'h14b7: char_row_bitmap <= 16'b0000000000000000;
		15'h14b8: char_row_bitmap <= 16'b0000000000000000;
		15'h14b9: char_row_bitmap <= 16'b0000000000000000;
		15'h14ba: char_row_bitmap <= 16'b0000000000000000;
		15'h14bb: char_row_bitmap <= 16'b0000000000000000;
		15'h14bc: char_row_bitmap <= 16'b0000000000000000;
		15'h14bd: char_row_bitmap <= 16'b0000000000000000;
		15'h14be: char_row_bitmap <= 16'b0000000000000000;
		15'h14bf: char_row_bitmap <= 16'b0000000000000000;
		15'h14c0: char_row_bitmap <= 16'b0000000000000000;
		15'h14c1: char_row_bitmap <= 16'b0000000000000000;
		15'h14c2: char_row_bitmap <= 16'b0000000000000000;
		15'h14c3: char_row_bitmap <= 16'b0000000000000000;
		15'h14c4: char_row_bitmap <= 16'b0000000000000000;
		15'h14c5: char_row_bitmap <= 16'b0000000000000000;
		15'h14c6: char_row_bitmap <= 16'b0000000000000000;
		15'h14c7: char_row_bitmap <= 16'b0000000000000000;
		15'h14c8: char_row_bitmap <= 16'b0000000000000000;
		15'h14c9: char_row_bitmap <= 16'b0000000000000000;
		15'h14ca: char_row_bitmap <= 16'b0000000000000000;
		15'h14cb: char_row_bitmap <= 16'b0000000000000000;
		15'h14cc: char_row_bitmap <= 16'b0000000000000000;
		15'h14cd: char_row_bitmap <= 16'b0000000000000000;
		15'h14ce: char_row_bitmap <= 16'b0000000000000000;
		15'h14cf: char_row_bitmap <= 16'b0000000000000000;
		15'h14d0: char_row_bitmap <= 16'b0000000000000000;
		15'h14d1: char_row_bitmap <= 16'b0000000000000000;
		15'h14d2: char_row_bitmap <= 16'b0000000000000000;
		15'h14d3: char_row_bitmap <= 16'b0000000000000000;
		15'h14d4: char_row_bitmap <= 16'b0000000000000000;
		15'h14d5: char_row_bitmap <= 16'b0000000000000000;
		15'h14d6: char_row_bitmap <= 16'b0000000000000000;
		15'h14d7: char_row_bitmap <= 16'b0000000000000000;
		15'h14d8: char_row_bitmap <= 16'b0000000000000000;
		15'h14d9: char_row_bitmap <= 16'b0000000000000000;
		15'h14da: char_row_bitmap <= 16'b0000000000000000;
		15'h14db: char_row_bitmap <= 16'b0000000000000000;
		15'h14dc: char_row_bitmap <= 16'b0000000000000000;
		15'h14dd: char_row_bitmap <= 16'b0000000000000000;
		15'h14de: char_row_bitmap <= 16'b0000000000000000;
		15'h14df: char_row_bitmap <= 16'b0000000000000000;
		15'h14e0: char_row_bitmap <= 16'b0000000000000000;
		15'h14e1: char_row_bitmap <= 16'b0000000000000000;
		15'h14e2: char_row_bitmap <= 16'b0000000000000000;
		15'h14e3: char_row_bitmap <= 16'b0000000000000000;
		15'h14e4: char_row_bitmap <= 16'b0000000000000000;
		15'h14e5: char_row_bitmap <= 16'b0000000000000000;
		15'h14e6: char_row_bitmap <= 16'b0000000000000000;
		15'h14e7: char_row_bitmap <= 16'b0000000000000000;
		15'h14e8: char_row_bitmap <= 16'b0000000000000000;
		15'h14e9: char_row_bitmap <= 16'b0000000000000000;
		15'h14ea: char_row_bitmap <= 16'b0000000000000000;
		15'h14eb: char_row_bitmap <= 16'b0000000000000000;
		15'h14ec: char_row_bitmap <= 16'b0000000000000000;
		15'h14ed: char_row_bitmap <= 16'b0000000000000000;
		15'h14ee: char_row_bitmap <= 16'b0000000000000000;
		15'h14ef: char_row_bitmap <= 16'b0000000000000000;
		15'h14f0: char_row_bitmap <= 16'b0000000000000000;
		15'h14f1: char_row_bitmap <= 16'b0000000000000000;
		15'h14f2: char_row_bitmap <= 16'b0000000000000000;
		15'h14f3: char_row_bitmap <= 16'b0000000000000000;
		15'h14f4: char_row_bitmap <= 16'b0000000000000000;
		15'h14f5: char_row_bitmap <= 16'b0000000000000000;
		15'h14f6: char_row_bitmap <= 16'b0000000000000000;
		15'h14f7: char_row_bitmap <= 16'b0000000000000000;
		15'h14f8: char_row_bitmap <= 16'b0000000000000000;
		15'h14f9: char_row_bitmap <= 16'b0000000000000000;
		15'h14fa: char_row_bitmap <= 16'b0000000000000000;
		15'h14fb: char_row_bitmap <= 16'b0000000000000000;
		15'h14fc: char_row_bitmap <= 16'b0000000000000000;
		15'h14fd: char_row_bitmap <= 16'b0000000000000000;
		15'h14fe: char_row_bitmap <= 16'b0000000000000000;
		15'h14ff: char_row_bitmap <= 16'b0000000000000000;
		15'h1500: char_row_bitmap <= 16'b0000000000000000;
		15'h1501: char_row_bitmap <= 16'b0000000000000000;
		15'h1502: char_row_bitmap <= 16'b0000000000000000;
		15'h1503: char_row_bitmap <= 16'b0000000000000000;
		15'h1504: char_row_bitmap <= 16'b0000000000000000;
		15'h1505: char_row_bitmap <= 16'b0000000000000000;
		15'h1506: char_row_bitmap <= 16'b0000000000000000;
		15'h1507: char_row_bitmap <= 16'b0000000000000000;
		15'h1508: char_row_bitmap <= 16'b0000000000000000;
		15'h1509: char_row_bitmap <= 16'b0000000000000000;
		15'h150a: char_row_bitmap <= 16'b0000000000000000;
		15'h150b: char_row_bitmap <= 16'b0000000000000000;
		15'h150c: char_row_bitmap <= 16'b0000000000000000;
		15'h150d: char_row_bitmap <= 16'b0000000000000000;
		15'h150e: char_row_bitmap <= 16'b0000000000000000;
		15'h150f: char_row_bitmap <= 16'b0000000000000000;
		15'h1510: char_row_bitmap <= 16'b0000000000000000;
		15'h1511: char_row_bitmap <= 16'b0000000000000000;
		15'h1512: char_row_bitmap <= 16'b0000000000000000;
		15'h1513: char_row_bitmap <= 16'b0000000000000000;
		15'h1514: char_row_bitmap <= 16'b0000000000000000;
		15'h1515: char_row_bitmap <= 16'b0000000000000000;
		15'h1516: char_row_bitmap <= 16'b0000000000000000;
		15'h1517: char_row_bitmap <= 16'b0000000000000000;
		15'h1518: char_row_bitmap <= 16'b0000000000000000;
		15'h1519: char_row_bitmap <= 16'b0000000000000000;
		15'h151a: char_row_bitmap <= 16'b0000000000000000;
		15'h151b: char_row_bitmap <= 16'b0000000000000000;
		15'h151c: char_row_bitmap <= 16'b0000000000000000;
		15'h151d: char_row_bitmap <= 16'b0000000000000000;
		15'h151e: char_row_bitmap <= 16'b0000000000000000;
		15'h151f: char_row_bitmap <= 16'b0000000000000000;
		15'h1520: char_row_bitmap <= 16'b0000000000000000;
		15'h1521: char_row_bitmap <= 16'b0000000000000000;
		15'h1522: char_row_bitmap <= 16'b0000000000000000;
		15'h1523: char_row_bitmap <= 16'b0000000000000000;
		15'h1524: char_row_bitmap <= 16'b0000000000000000;
		15'h1525: char_row_bitmap <= 16'b0000000000000000;
		15'h1526: char_row_bitmap <= 16'b0000000000000000;
		15'h1527: char_row_bitmap <= 16'b0000000000000000;
		15'h1528: char_row_bitmap <= 16'b0000000000000000;
		15'h1529: char_row_bitmap <= 16'b0000000000000000;
		15'h152a: char_row_bitmap <= 16'b0000000000000000;
		15'h152b: char_row_bitmap <= 16'b0000000000000000;
		15'h152c: char_row_bitmap <= 16'b0000000000000000;
		15'h152d: char_row_bitmap <= 16'b0000000000000000;
		15'h152e: char_row_bitmap <= 16'b0000000000000000;
		15'h152f: char_row_bitmap <= 16'b0000000000000000;
		15'h1530: char_row_bitmap <= 16'b0000000000000000;
		15'h1531: char_row_bitmap <= 16'b0000000000000000;
		15'h1532: char_row_bitmap <= 16'b0000000000000000;
		15'h1533: char_row_bitmap <= 16'b0000000000000000;
		15'h1534: char_row_bitmap <= 16'b0000000000000000;
		15'h1535: char_row_bitmap <= 16'b0000000000000000;
		15'h1536: char_row_bitmap <= 16'b0000000000000000;
		15'h1537: char_row_bitmap <= 16'b0000000000000000;
		15'h1538: char_row_bitmap <= 16'b0000000000000000;
		15'h1539: char_row_bitmap <= 16'b0000000000000000;
		15'h153a: char_row_bitmap <= 16'b0000000000000000;
		15'h153b: char_row_bitmap <= 16'b0000000000000000;
		15'h153c: char_row_bitmap <= 16'b0000000000000000;
		15'h153d: char_row_bitmap <= 16'b0000000000000000;
		15'h153e: char_row_bitmap <= 16'b0000000000000000;
		15'h153f: char_row_bitmap <= 16'b0000000000000000;
		15'h1540: char_row_bitmap <= 16'b0000000000000000;
		15'h1541: char_row_bitmap <= 16'b0000000000000000;
		15'h1542: char_row_bitmap <= 16'b0000000000000000;
		15'h1543: char_row_bitmap <= 16'b0000000000000000;
		15'h1544: char_row_bitmap <= 16'b0000000000000000;
		15'h1545: char_row_bitmap <= 16'b0000000000000000;
		15'h1546: char_row_bitmap <= 16'b0000000000000000;
		15'h1547: char_row_bitmap <= 16'b0000000000000000;
		15'h1548: char_row_bitmap <= 16'b0000000000000000;
		15'h1549: char_row_bitmap <= 16'b0000000000000000;
		15'h154a: char_row_bitmap <= 16'b0000000000000000;
		15'h154b: char_row_bitmap <= 16'b0000000000000000;
		15'h154c: char_row_bitmap <= 16'b0000000000000000;
		15'h154d: char_row_bitmap <= 16'b0000000000000000;
		15'h154e: char_row_bitmap <= 16'b0000000000000000;
		15'h154f: char_row_bitmap <= 16'b0000000000000000;
		15'h1550: char_row_bitmap <= 16'b0000000000000000;
		15'h1551: char_row_bitmap <= 16'b0000000000000000;
		15'h1552: char_row_bitmap <= 16'b0000000000000000;
		15'h1553: char_row_bitmap <= 16'b0000000000000000;
		15'h1554: char_row_bitmap <= 16'b0000000000000000;
		15'h1555: char_row_bitmap <= 16'b0000000000000000;
		15'h1556: char_row_bitmap <= 16'b0000000000000000;
		15'h1557: char_row_bitmap <= 16'b0000000000000000;
		15'h1558: char_row_bitmap <= 16'b0000000000000000;
		15'h1559: char_row_bitmap <= 16'b0000000000000000;
		15'h155a: char_row_bitmap <= 16'b0000000000000000;
		15'h155b: char_row_bitmap <= 16'b0000000000000000;
		15'h155c: char_row_bitmap <= 16'b0000000000000000;
		15'h155d: char_row_bitmap <= 16'b0000000000000000;
		15'h155e: char_row_bitmap <= 16'b0000000000000000;
		15'h155f: char_row_bitmap <= 16'b0000000000000000;
		15'h1560: char_row_bitmap <= 16'b0000000000000000;
		15'h1561: char_row_bitmap <= 16'b0000000000000000;
		15'h1562: char_row_bitmap <= 16'b0000000000000000;
		15'h1563: char_row_bitmap <= 16'b0000000000000000;
		15'h1564: char_row_bitmap <= 16'b0000000000000000;
		15'h1565: char_row_bitmap <= 16'b0000000000000000;
		15'h1566: char_row_bitmap <= 16'b0000000000000000;
		15'h1567: char_row_bitmap <= 16'b0000000000000000;
		15'h1568: char_row_bitmap <= 16'b0000000000000000;
		15'h1569: char_row_bitmap <= 16'b0000000000000000;
		15'h156a: char_row_bitmap <= 16'b0000000000000000;
		15'h156b: char_row_bitmap <= 16'b0000000000000000;
		15'h156c: char_row_bitmap <= 16'b0000000000000000;
		15'h156d: char_row_bitmap <= 16'b0000000000000000;
		15'h156e: char_row_bitmap <= 16'b0000000000000000;
		15'h156f: char_row_bitmap <= 16'b0000000000000000;
		15'h1570: char_row_bitmap <= 16'b0000000000000000;
		15'h1571: char_row_bitmap <= 16'b0000000000000000;
		15'h1572: char_row_bitmap <= 16'b0000000000000000;
		15'h1573: char_row_bitmap <= 16'b0000000000000000;
		15'h1574: char_row_bitmap <= 16'b0000000000000000;
		15'h1575: char_row_bitmap <= 16'b0000000000000000;
		15'h1576: char_row_bitmap <= 16'b0000000000000000;
		15'h1577: char_row_bitmap <= 16'b0000000000000000;
		15'h1578: char_row_bitmap <= 16'b0000000000000000;
		15'h1579: char_row_bitmap <= 16'b0000000000000000;
		15'h157a: char_row_bitmap <= 16'b0000000000000000;
		15'h157b: char_row_bitmap <= 16'b0000000000000000;
		15'h157c: char_row_bitmap <= 16'b0000000000000000;
		15'h157d: char_row_bitmap <= 16'b0000000000000000;
		15'h157e: char_row_bitmap <= 16'b0000000000000000;
		15'h157f: char_row_bitmap <= 16'b0000000000000000;
		15'h1580: char_row_bitmap <= 16'b0000000000000000;
		15'h1581: char_row_bitmap <= 16'b0000000000000000;
		15'h1582: char_row_bitmap <= 16'b0000000000000000;
		15'h1583: char_row_bitmap <= 16'b0000000000000000;
		15'h1584: char_row_bitmap <= 16'b0000000000000000;
		15'h1585: char_row_bitmap <= 16'b0000000000000000;
		15'h1586: char_row_bitmap <= 16'b0000000000000000;
		15'h1587: char_row_bitmap <= 16'b0000000000000000;
		15'h1588: char_row_bitmap <= 16'b0000000000000000;
		15'h1589: char_row_bitmap <= 16'b0000000000000000;
		15'h158a: char_row_bitmap <= 16'b0000000000000000;
		15'h158b: char_row_bitmap <= 16'b0000000000000000;
		15'h158c: char_row_bitmap <= 16'b0000000000000000;
		15'h158d: char_row_bitmap <= 16'b0000000000000000;
		15'h158e: char_row_bitmap <= 16'b0000000000000000;
		15'h158f: char_row_bitmap <= 16'b0000000000000000;
		15'h1590: char_row_bitmap <= 16'b0000000000000000;
		15'h1591: char_row_bitmap <= 16'b0000000000000000;
		15'h1592: char_row_bitmap <= 16'b0000000000000000;
		15'h1593: char_row_bitmap <= 16'b0000000000000000;
		15'h1594: char_row_bitmap <= 16'b0000000000000000;
		15'h1595: char_row_bitmap <= 16'b0000000000000000;
		15'h1596: char_row_bitmap <= 16'b0000000000000000;
		15'h1597: char_row_bitmap <= 16'b0000000000000000;
		15'h1598: char_row_bitmap <= 16'b0000000000000000;
		15'h1599: char_row_bitmap <= 16'b0000000000000000;
		15'h159a: char_row_bitmap <= 16'b0000000000000000;
		15'h159b: char_row_bitmap <= 16'b0000000000000000;
		15'h159c: char_row_bitmap <= 16'b0000000000000000;
		15'h159d: char_row_bitmap <= 16'b0000000000000000;
		15'h159e: char_row_bitmap <= 16'b0000000000000000;
		15'h159f: char_row_bitmap <= 16'b0000000000000000;
		15'h15a0: char_row_bitmap <= 16'b0000000000000000;
		15'h15a1: char_row_bitmap <= 16'b0000000000000000;
		15'h15a2: char_row_bitmap <= 16'b0000000000000000;
		15'h15a3: char_row_bitmap <= 16'b0000000000000000;
		15'h15a4: char_row_bitmap <= 16'b0000000000000000;
		15'h15a5: char_row_bitmap <= 16'b0000000000000000;
		15'h15a6: char_row_bitmap <= 16'b0000000000000000;
		15'h15a7: char_row_bitmap <= 16'b0000000000000000;
		15'h15a8: char_row_bitmap <= 16'b0000000000000000;
		15'h15a9: char_row_bitmap <= 16'b0000000000000000;
		15'h15aa: char_row_bitmap <= 16'b0000000000000000;
		15'h15ab: char_row_bitmap <= 16'b0000000000000000;
		15'h15ac: char_row_bitmap <= 16'b0000000000000000;
		15'h15ad: char_row_bitmap <= 16'b0000000000000000;
		15'h15ae: char_row_bitmap <= 16'b0000000000000000;
		15'h15af: char_row_bitmap <= 16'b0000000000000000;
		15'h15b0: char_row_bitmap <= 16'b0000000000000000;
		15'h15b1: char_row_bitmap <= 16'b0000000000000000;
		15'h15b2: char_row_bitmap <= 16'b0000000000000000;
		15'h15b3: char_row_bitmap <= 16'b0000000000000000;
		15'h15b4: char_row_bitmap <= 16'b0000000000000000;
		15'h15b5: char_row_bitmap <= 16'b0000000000000000;
		15'h15b6: char_row_bitmap <= 16'b0000000000000000;
		15'h15b7: char_row_bitmap <= 16'b0000000000000000;
		15'h15b8: char_row_bitmap <= 16'b0000000000000000;
		15'h15b9: char_row_bitmap <= 16'b0000000000000000;
		15'h15ba: char_row_bitmap <= 16'b0000000000000000;
		15'h15bb: char_row_bitmap <= 16'b0000000000000000;
		15'h15bc: char_row_bitmap <= 16'b0000000000000000;
		15'h15bd: char_row_bitmap <= 16'b0000000000000000;
		15'h15be: char_row_bitmap <= 16'b0000000000000000;
		15'h15bf: char_row_bitmap <= 16'b0000000000000000;
		15'h15c0: char_row_bitmap <= 16'b0000000000000000;
		15'h15c1: char_row_bitmap <= 16'b0000000000000000;
		15'h15c2: char_row_bitmap <= 16'b0000000000000000;
		15'h15c3: char_row_bitmap <= 16'b0000000000000000;
		15'h15c4: char_row_bitmap <= 16'b0000000000000000;
		15'h15c5: char_row_bitmap <= 16'b0000000000000000;
		15'h15c6: char_row_bitmap <= 16'b0000000000000000;
		15'h15c7: char_row_bitmap <= 16'b0000000000000000;
		15'h15c8: char_row_bitmap <= 16'b0000000000000000;
		15'h15c9: char_row_bitmap <= 16'b0000000000000000;
		15'h15ca: char_row_bitmap <= 16'b0000000000000000;
		15'h15cb: char_row_bitmap <= 16'b0000000000000000;
		15'h15cc: char_row_bitmap <= 16'b0000000000000000;
		15'h15cd: char_row_bitmap <= 16'b0000000000000000;
		15'h15ce: char_row_bitmap <= 16'b0000000000000000;
		15'h15cf: char_row_bitmap <= 16'b0000000000000000;
		15'h15d0: char_row_bitmap <= 16'b0000000000000000;
		15'h15d1: char_row_bitmap <= 16'b0000000000000000;
		15'h15d2: char_row_bitmap <= 16'b0000000000000000;
		15'h15d3: char_row_bitmap <= 16'b0000000000000000;
		15'h15d4: char_row_bitmap <= 16'b0000000000000000;
		15'h15d5: char_row_bitmap <= 16'b0000000000000000;
		15'h15d6: char_row_bitmap <= 16'b0000000000000000;
		15'h15d7: char_row_bitmap <= 16'b0000000000000000;
		15'h15d8: char_row_bitmap <= 16'b0000000000000000;
		15'h15d9: char_row_bitmap <= 16'b0000000000000000;
		15'h15da: char_row_bitmap <= 16'b0000000000000000;
		15'h15db: char_row_bitmap <= 16'b0000000000000000;
		15'h15dc: char_row_bitmap <= 16'b0000000000000000;
		15'h15dd: char_row_bitmap <= 16'b0000000000000000;
		15'h15de: char_row_bitmap <= 16'b0000000000000000;
		15'h15df: char_row_bitmap <= 16'b0000000000000000;
		15'h15e0: char_row_bitmap <= 16'b0000000000000000;
		15'h15e1: char_row_bitmap <= 16'b0000000000000000;
		15'h15e2: char_row_bitmap <= 16'b0000000000000000;
		15'h15e3: char_row_bitmap <= 16'b0000000000000000;
		15'h15e4: char_row_bitmap <= 16'b0000000000000000;
		15'h15e5: char_row_bitmap <= 16'b0000000000000000;
		15'h15e6: char_row_bitmap <= 16'b0000000000000000;
		15'h15e7: char_row_bitmap <= 16'b0000000000000000;
		15'h15e8: char_row_bitmap <= 16'b0000000000000000;
		15'h15e9: char_row_bitmap <= 16'b0000000000000000;
		15'h15ea: char_row_bitmap <= 16'b0000000000000000;
		15'h15eb: char_row_bitmap <= 16'b0000000000000000;
		15'h15ec: char_row_bitmap <= 16'b0000000000000000;
		15'h15ed: char_row_bitmap <= 16'b0000000000000000;
		15'h15ee: char_row_bitmap <= 16'b0000000000000000;
		15'h15ef: char_row_bitmap <= 16'b0000000000000000;
		15'h15f0: char_row_bitmap <= 16'b0000000000000000;
		15'h15f1: char_row_bitmap <= 16'b0000000000000000;
		15'h15f2: char_row_bitmap <= 16'b0000000000000000;
		15'h15f3: char_row_bitmap <= 16'b0000000000000000;
		15'h15f4: char_row_bitmap <= 16'b0000000000000000;
		15'h15f5: char_row_bitmap <= 16'b0000000000000000;
		15'h15f6: char_row_bitmap <= 16'b0000000000000000;
		15'h15f7: char_row_bitmap <= 16'b0000000000000000;
		15'h15f8: char_row_bitmap <= 16'b0000000000000000;
		15'h15f9: char_row_bitmap <= 16'b0000000000000000;
		15'h15fa: char_row_bitmap <= 16'b0000000000000000;
		15'h15fb: char_row_bitmap <= 16'b0000000000000000;
		15'h15fc: char_row_bitmap <= 16'b0000000000000000;
		15'h15fd: char_row_bitmap <= 16'b0000000000000000;
		15'h15fe: char_row_bitmap <= 16'b0000000000000000;
		15'h15ff: char_row_bitmap <= 16'b0000000000000000;
		15'h1600: char_row_bitmap <= 16'b0000000000000000;
		15'h1601: char_row_bitmap <= 16'b0000000000000000;
		15'h1602: char_row_bitmap <= 16'b0000000000000000;
		15'h1603: char_row_bitmap <= 16'b0000000000000000;
		15'h1604: char_row_bitmap <= 16'b0000000000000000;
		15'h1605: char_row_bitmap <= 16'b0000000000000000;
		15'h1606: char_row_bitmap <= 16'b0000000000000000;
		15'h1607: char_row_bitmap <= 16'b0000000000000000;
		15'h1608: char_row_bitmap <= 16'b0000000000000000;
		15'h1609: char_row_bitmap <= 16'b0000000000000000;
		15'h160a: char_row_bitmap <= 16'b0000000000000000;
		15'h160b: char_row_bitmap <= 16'b0000000000000000;
		15'h160c: char_row_bitmap <= 16'b0000000000000000;
		15'h160d: char_row_bitmap <= 16'b0000000000000000;
		15'h160e: char_row_bitmap <= 16'b0000000000000000;
		15'h160f: char_row_bitmap <= 16'b0000000000000000;
		15'h1610: char_row_bitmap <= 16'b0000000000000000;
		15'h1611: char_row_bitmap <= 16'b0000000000000000;
		15'h1612: char_row_bitmap <= 16'b0000000000000000;
		15'h1613: char_row_bitmap <= 16'b0000000000000000;
		15'h1614: char_row_bitmap <= 16'b0000000000000000;
		15'h1615: char_row_bitmap <= 16'b0000000000000000;
		15'h1616: char_row_bitmap <= 16'b0000000000000000;
		15'h1617: char_row_bitmap <= 16'b0000000000000000;
		15'h1618: char_row_bitmap <= 16'b0000000000000000;
		15'h1619: char_row_bitmap <= 16'b0000000000000000;
		15'h161a: char_row_bitmap <= 16'b0000000000000000;
		15'h161b: char_row_bitmap <= 16'b0000000000000000;
		15'h161c: char_row_bitmap <= 16'b0000000000000000;
		15'h161d: char_row_bitmap <= 16'b0000000000000000;
		15'h161e: char_row_bitmap <= 16'b0000000000000000;
		15'h161f: char_row_bitmap <= 16'b0000000000000000;
		15'h1620: char_row_bitmap <= 16'b0000000000000000;
		15'h1621: char_row_bitmap <= 16'b0000000000000000;
		15'h1622: char_row_bitmap <= 16'b0000000000000000;
		15'h1623: char_row_bitmap <= 16'b0000000000000000;
		15'h1624: char_row_bitmap <= 16'b0000000000000000;
		15'h1625: char_row_bitmap <= 16'b0000000000000000;
		15'h1626: char_row_bitmap <= 16'b0000000000000000;
		15'h1627: char_row_bitmap <= 16'b0000000000000000;
		15'h1628: char_row_bitmap <= 16'b0000000000000000;
		15'h1629: char_row_bitmap <= 16'b0000000000000000;
		15'h162a: char_row_bitmap <= 16'b0000000000000000;
		15'h162b: char_row_bitmap <= 16'b0000000000000000;
		15'h162c: char_row_bitmap <= 16'b0000000000000000;
		15'h162d: char_row_bitmap <= 16'b0000000000000000;
		15'h162e: char_row_bitmap <= 16'b0000000000000000;
		15'h162f: char_row_bitmap <= 16'b0000000000000000;
		15'h1630: char_row_bitmap <= 16'b0000000000000000;
		15'h1631: char_row_bitmap <= 16'b0000000000000000;
		15'h1632: char_row_bitmap <= 16'b0000000000000000;
		15'h1633: char_row_bitmap <= 16'b0000000000000000;
		15'h1634: char_row_bitmap <= 16'b0000000000000000;
		15'h1635: char_row_bitmap <= 16'b0000000000000000;
		15'h1636: char_row_bitmap <= 16'b0000000000000000;
		15'h1637: char_row_bitmap <= 16'b0000000000000000;
		15'h1638: char_row_bitmap <= 16'b0000000000000000;
		15'h1639: char_row_bitmap <= 16'b0000000000000000;
		15'h163a: char_row_bitmap <= 16'b0000000000000000;
		15'h163b: char_row_bitmap <= 16'b0000000000000000;
		15'h163c: char_row_bitmap <= 16'b0000000000000000;
		15'h163d: char_row_bitmap <= 16'b0000000000000000;
		15'h163e: char_row_bitmap <= 16'b0000000000000000;
		15'h163f: char_row_bitmap <= 16'b0000000000000000;
		15'h1640: char_row_bitmap <= 16'b0000000000000000;
		15'h1641: char_row_bitmap <= 16'b0000000000000000;
		15'h1642: char_row_bitmap <= 16'b0000000000000000;
		15'h1643: char_row_bitmap <= 16'b0000000000000000;
		15'h1644: char_row_bitmap <= 16'b0000000000000000;
		15'h1645: char_row_bitmap <= 16'b0000000000000000;
		15'h1646: char_row_bitmap <= 16'b0000000000000000;
		15'h1647: char_row_bitmap <= 16'b0000000000000000;
		15'h1648: char_row_bitmap <= 16'b0000000000000000;
		15'h1649: char_row_bitmap <= 16'b0000000000000000;
		15'h164a: char_row_bitmap <= 16'b0000000000000000;
		15'h164b: char_row_bitmap <= 16'b0000000000000000;
		15'h164c: char_row_bitmap <= 16'b0000000000000000;
		15'h164d: char_row_bitmap <= 16'b0000000000000000;
		15'h164e: char_row_bitmap <= 16'b0000000000000000;
		15'h164f: char_row_bitmap <= 16'b0000000000000000;
		15'h1650: char_row_bitmap <= 16'b0000000000000000;
		15'h1651: char_row_bitmap <= 16'b0000000000000000;
		15'h1652: char_row_bitmap <= 16'b0000000000000000;
		15'h1653: char_row_bitmap <= 16'b0000000000000000;
		15'h1654: char_row_bitmap <= 16'b0000000000000000;
		15'h1655: char_row_bitmap <= 16'b0000000000000000;
		15'h1656: char_row_bitmap <= 16'b0000000000000000;
		15'h1657: char_row_bitmap <= 16'b0000000000000000;
		15'h1658: char_row_bitmap <= 16'b0000000000000000;
		15'h1659: char_row_bitmap <= 16'b0000000000000000;
		15'h165a: char_row_bitmap <= 16'b0000000000000000;
		15'h165b: char_row_bitmap <= 16'b0000000000000000;
		15'h165c: char_row_bitmap <= 16'b0000000000000000;
		15'h165d: char_row_bitmap <= 16'b0000000000000000;
		15'h165e: char_row_bitmap <= 16'b0000000000000000;
		15'h165f: char_row_bitmap <= 16'b0000000000000000;
		15'h1660: char_row_bitmap <= 16'b0000000000000000;
		15'h1661: char_row_bitmap <= 16'b0000000000000000;
		15'h1662: char_row_bitmap <= 16'b0000000000000000;
		15'h1663: char_row_bitmap <= 16'b0000000000000000;
		15'h1664: char_row_bitmap <= 16'b0000000000000000;
		15'h1665: char_row_bitmap <= 16'b0000000000000000;
		15'h1666: char_row_bitmap <= 16'b0000000000000000;
		15'h1667: char_row_bitmap <= 16'b0000000000000000;
		15'h1668: char_row_bitmap <= 16'b0000000000000000;
		15'h1669: char_row_bitmap <= 16'b0000000000000000;
		15'h166a: char_row_bitmap <= 16'b0000000000000000;
		15'h166b: char_row_bitmap <= 16'b0000000000000000;
		15'h166c: char_row_bitmap <= 16'b0000000000000000;
		15'h166d: char_row_bitmap <= 16'b0000000000000000;
		15'h166e: char_row_bitmap <= 16'b0000000000000000;
		15'h166f: char_row_bitmap <= 16'b0000000000000000;
		15'h1670: char_row_bitmap <= 16'b0000000000000000;
		15'h1671: char_row_bitmap <= 16'b0000000000000000;
		15'h1672: char_row_bitmap <= 16'b0000000000000000;
		15'h1673: char_row_bitmap <= 16'b0000000000000000;
		15'h1674: char_row_bitmap <= 16'b0000000000000000;
		15'h1675: char_row_bitmap <= 16'b0000000000000000;
		15'h1676: char_row_bitmap <= 16'b0000000000000000;
		15'h1677: char_row_bitmap <= 16'b0000000000000000;
		15'h1678: char_row_bitmap <= 16'b0000000000000000;
		15'h1679: char_row_bitmap <= 16'b0000000000000000;
		15'h167a: char_row_bitmap <= 16'b0000000000000000;
		15'h167b: char_row_bitmap <= 16'b0000000000000000;
		15'h167c: char_row_bitmap <= 16'b0000000000000000;
		15'h167d: char_row_bitmap <= 16'b0000000000000000;
		15'h167e: char_row_bitmap <= 16'b0000000000000000;
		15'h167f: char_row_bitmap <= 16'b0000000000000000;
		15'h1680: char_row_bitmap <= 16'b0000000000000000;
		15'h1681: char_row_bitmap <= 16'b0000000000000000;
		15'h1682: char_row_bitmap <= 16'b0000000000000000;
		15'h1683: char_row_bitmap <= 16'b0000000000000000;
		15'h1684: char_row_bitmap <= 16'b0000000000000000;
		15'h1685: char_row_bitmap <= 16'b0000000000000000;
		15'h1686: char_row_bitmap <= 16'b0000000000000000;
		15'h1687: char_row_bitmap <= 16'b0000000000000000;
		15'h1688: char_row_bitmap <= 16'b0000000000000000;
		15'h1689: char_row_bitmap <= 16'b0000000000000000;
		15'h168a: char_row_bitmap <= 16'b0000000000000000;
		15'h168b: char_row_bitmap <= 16'b0000000000000000;
		15'h168c: char_row_bitmap <= 16'b0000000000000000;
		15'h168d: char_row_bitmap <= 16'b0000000000000000;
		15'h168e: char_row_bitmap <= 16'b0000000000000000;
		15'h168f: char_row_bitmap <= 16'b0000000000000000;
		15'h1690: char_row_bitmap <= 16'b0000000000000000;
		15'h1691: char_row_bitmap <= 16'b0000000000000000;
		15'h1692: char_row_bitmap <= 16'b0000000000000000;
		15'h1693: char_row_bitmap <= 16'b0000000000000000;
		15'h1694: char_row_bitmap <= 16'b0000000000000000;
		15'h1695: char_row_bitmap <= 16'b0000000000000000;
		15'h1696: char_row_bitmap <= 16'b0000000000000000;
		15'h1697: char_row_bitmap <= 16'b0000000000000000;
		15'h1698: char_row_bitmap <= 16'b0000000000000000;
		15'h1699: char_row_bitmap <= 16'b0000000000000000;
		15'h169a: char_row_bitmap <= 16'b0000000000000000;
		15'h169b: char_row_bitmap <= 16'b0000000000000000;
		15'h169c: char_row_bitmap <= 16'b0000000000000000;
		15'h169d: char_row_bitmap <= 16'b0000000000000000;
		15'h169e: char_row_bitmap <= 16'b0000000000000000;
		15'h169f: char_row_bitmap <= 16'b0000000000000000;
		15'h16a0: char_row_bitmap <= 16'b0000000000000000;
		15'h16a1: char_row_bitmap <= 16'b0000000000000000;
		15'h16a2: char_row_bitmap <= 16'b0000000000000000;
		15'h16a3: char_row_bitmap <= 16'b0000000000000000;
		15'h16a4: char_row_bitmap <= 16'b0000000000000000;
		15'h16a5: char_row_bitmap <= 16'b0000000000000000;
		15'h16a6: char_row_bitmap <= 16'b0000000000000000;
		15'h16a7: char_row_bitmap <= 16'b0000000000000000;
		15'h16a8: char_row_bitmap <= 16'b0000000000000000;
		15'h16a9: char_row_bitmap <= 16'b0000000000000000;
		15'h16aa: char_row_bitmap <= 16'b0000000000000000;
		15'h16ab: char_row_bitmap <= 16'b0000000000000000;
		15'h16ac: char_row_bitmap <= 16'b0000000000000000;
		15'h16ad: char_row_bitmap <= 16'b0000000000000000;
		15'h16ae: char_row_bitmap <= 16'b0000000000000000;
		15'h16af: char_row_bitmap <= 16'b0000000000000000;
		15'h16b0: char_row_bitmap <= 16'b0000000000000000;
		15'h16b1: char_row_bitmap <= 16'b0000000000000000;
		15'h16b2: char_row_bitmap <= 16'b0000000000000000;
		15'h16b3: char_row_bitmap <= 16'b0000000000000000;
		15'h16b4: char_row_bitmap <= 16'b0000000000000000;
		15'h16b5: char_row_bitmap <= 16'b0000000000000000;
		15'h16b6: char_row_bitmap <= 16'b0000000000000000;
		15'h16b7: char_row_bitmap <= 16'b0000000000000000;
		15'h16b8: char_row_bitmap <= 16'b0000000000000000;
		15'h16b9: char_row_bitmap <= 16'b0000000000000000;
		15'h16ba: char_row_bitmap <= 16'b0000000000000000;
		15'h16bb: char_row_bitmap <= 16'b0000000000000000;
		15'h16bc: char_row_bitmap <= 16'b0000000000000000;
		15'h16bd: char_row_bitmap <= 16'b0000000000000000;
		15'h16be: char_row_bitmap <= 16'b0000000000000000;
		15'h16bf: char_row_bitmap <= 16'b0000000000000000;
		15'h16c0: char_row_bitmap <= 16'b0000000000000000;
		15'h16c1: char_row_bitmap <= 16'b0000000000000000;
		15'h16c2: char_row_bitmap <= 16'b0000000000000000;
		15'h16c3: char_row_bitmap <= 16'b0000000000000000;
		15'h16c4: char_row_bitmap <= 16'b0000000000000000;
		15'h16c5: char_row_bitmap <= 16'b0000000000000000;
		15'h16c6: char_row_bitmap <= 16'b0000000000000000;
		15'h16c7: char_row_bitmap <= 16'b0000000000000000;
		15'h16c8: char_row_bitmap <= 16'b0000000000000000;
		15'h16c9: char_row_bitmap <= 16'b0000000000000000;
		15'h16ca: char_row_bitmap <= 16'b0000000000000000;
		15'h16cb: char_row_bitmap <= 16'b0000000000000000;
		15'h16cc: char_row_bitmap <= 16'b0000000000000000;
		15'h16cd: char_row_bitmap <= 16'b0000000000000000;
		15'h16ce: char_row_bitmap <= 16'b0000000000000000;
		15'h16cf: char_row_bitmap <= 16'b0000000000000000;
		15'h16d0: char_row_bitmap <= 16'b0000000000000000;
		15'h16d1: char_row_bitmap <= 16'b0000000000000000;
		15'h16d2: char_row_bitmap <= 16'b0000000000000000;
		15'h16d3: char_row_bitmap <= 16'b0000000000000000;
		15'h16d4: char_row_bitmap <= 16'b0000000000000000;
		15'h16d5: char_row_bitmap <= 16'b0000000000000000;
		15'h16d6: char_row_bitmap <= 16'b0000000000000000;
		15'h16d7: char_row_bitmap <= 16'b0000000000000000;
		15'h16d8: char_row_bitmap <= 16'b0000000000000000;
		15'h16d9: char_row_bitmap <= 16'b0000000000000000;
		15'h16da: char_row_bitmap <= 16'b0000000000000000;
		15'h16db: char_row_bitmap <= 16'b0000000000000000;
		15'h16dc: char_row_bitmap <= 16'b0000000000000000;
		15'h16dd: char_row_bitmap <= 16'b0000000000000000;
		15'h16de: char_row_bitmap <= 16'b0000000000000000;
		15'h16df: char_row_bitmap <= 16'b0000000000000000;
		15'h16e0: char_row_bitmap <= 16'b0000000000000000;
		15'h16e1: char_row_bitmap <= 16'b0000000000000000;
		15'h16e2: char_row_bitmap <= 16'b0000000000000000;
		15'h16e3: char_row_bitmap <= 16'b0000000000000000;
		15'h16e4: char_row_bitmap <= 16'b0000000000000000;
		15'h16e5: char_row_bitmap <= 16'b0000000000000000;
		15'h16e6: char_row_bitmap <= 16'b0000000000000000;
		15'h16e7: char_row_bitmap <= 16'b0000000000000000;
		15'h16e8: char_row_bitmap <= 16'b0000000000000000;
		15'h16e9: char_row_bitmap <= 16'b0000000000000000;
		15'h16ea: char_row_bitmap <= 16'b0000000000000000;
		15'h16eb: char_row_bitmap <= 16'b0000000000000000;
		15'h16ec: char_row_bitmap <= 16'b0000000000000000;
		15'h16ed: char_row_bitmap <= 16'b0000000000000000;
		15'h16ee: char_row_bitmap <= 16'b0000000000000000;
		15'h16ef: char_row_bitmap <= 16'b0000000000000000;
		15'h16f0: char_row_bitmap <= 16'b0000000000000000;
		15'h16f1: char_row_bitmap <= 16'b0000000000000000;
		15'h16f2: char_row_bitmap <= 16'b0000000000000000;
		15'h16f3: char_row_bitmap <= 16'b0000000000000000;
		15'h16f4: char_row_bitmap <= 16'b0000000000000000;
		15'h16f5: char_row_bitmap <= 16'b0000000000000000;
		15'h16f6: char_row_bitmap <= 16'b0000000000000000;
		15'h16f7: char_row_bitmap <= 16'b0000000000000000;
		15'h16f8: char_row_bitmap <= 16'b0000000000000000;
		15'h16f9: char_row_bitmap <= 16'b0000000000000000;
		15'h16fa: char_row_bitmap <= 16'b0000000000000000;
		15'h16fb: char_row_bitmap <= 16'b0000000000000000;
		15'h16fc: char_row_bitmap <= 16'b0000000000000000;
		15'h16fd: char_row_bitmap <= 16'b0000000000000000;
		15'h16fe: char_row_bitmap <= 16'b0000000000000000;
		15'h16ff: char_row_bitmap <= 16'b0000000000000000;
		15'h1700: char_row_bitmap <= 16'b0000000000000000;
		15'h1701: char_row_bitmap <= 16'b0000000000000000;
		15'h1702: char_row_bitmap <= 16'b0000000000000000;
		15'h1703: char_row_bitmap <= 16'b0000000000000000;
		15'h1704: char_row_bitmap <= 16'b0000000000000000;
		15'h1705: char_row_bitmap <= 16'b0000000000000000;
		15'h1706: char_row_bitmap <= 16'b0000000000000000;
		15'h1707: char_row_bitmap <= 16'b0000000000000000;
		15'h1708: char_row_bitmap <= 16'b0000000000000000;
		15'h1709: char_row_bitmap <= 16'b0000000000000000;
		15'h170a: char_row_bitmap <= 16'b0000000000000000;
		15'h170b: char_row_bitmap <= 16'b0000000000000000;
		15'h170c: char_row_bitmap <= 16'b0000000000000000;
		15'h170d: char_row_bitmap <= 16'b0000000000000000;
		15'h170e: char_row_bitmap <= 16'b0000000000000000;
		15'h170f: char_row_bitmap <= 16'b0000000000000000;
		15'h1710: char_row_bitmap <= 16'b0000000000000000;
		15'h1711: char_row_bitmap <= 16'b0000000000000000;
		15'h1712: char_row_bitmap <= 16'b0000000000000000;
		15'h1713: char_row_bitmap <= 16'b0000000000000000;
		15'h1714: char_row_bitmap <= 16'b0000000000000000;
		15'h1715: char_row_bitmap <= 16'b0000000000000000;
		15'h1716: char_row_bitmap <= 16'b0000000000000000;
		15'h1717: char_row_bitmap <= 16'b0000000000000000;
		15'h1718: char_row_bitmap <= 16'b0000000000000000;
		15'h1719: char_row_bitmap <= 16'b0000000000000000;
		15'h171a: char_row_bitmap <= 16'b0000000000000000;
		15'h171b: char_row_bitmap <= 16'b0000000000000000;
		15'h171c: char_row_bitmap <= 16'b0000000000000000;
		15'h171d: char_row_bitmap <= 16'b0000000000000000;
		15'h171e: char_row_bitmap <= 16'b0000000000000000;
		15'h171f: char_row_bitmap <= 16'b0000000000000000;
		15'h1720: char_row_bitmap <= 16'b0000000000000000;
		15'h1721: char_row_bitmap <= 16'b0000000000000000;
		15'h1722: char_row_bitmap <= 16'b0000000000000000;
		15'h1723: char_row_bitmap <= 16'b0000000000000000;
		15'h1724: char_row_bitmap <= 16'b0000000000000000;
		15'h1725: char_row_bitmap <= 16'b0000000000000000;
		15'h1726: char_row_bitmap <= 16'b0000000000000000;
		15'h1727: char_row_bitmap <= 16'b0000000000000000;
		15'h1728: char_row_bitmap <= 16'b0000000000000000;
		15'h1729: char_row_bitmap <= 16'b0000000000000000;
		15'h172a: char_row_bitmap <= 16'b0000000000000000;
		15'h172b: char_row_bitmap <= 16'b0000000000000000;
		15'h172c: char_row_bitmap <= 16'b0000000000000000;
		15'h172d: char_row_bitmap <= 16'b0000000000000000;
		15'h172e: char_row_bitmap <= 16'b0000000000000000;
		15'h172f: char_row_bitmap <= 16'b0000000000000000;
		15'h1730: char_row_bitmap <= 16'b0000000000000000;
		15'h1731: char_row_bitmap <= 16'b0000000000000000;
		15'h1732: char_row_bitmap <= 16'b0000000000000000;
		15'h1733: char_row_bitmap <= 16'b0000000000000000;
		15'h1734: char_row_bitmap <= 16'b0000000000000000;
		15'h1735: char_row_bitmap <= 16'b0000000000000000;
		15'h1736: char_row_bitmap <= 16'b0000000000000000;
		15'h1737: char_row_bitmap <= 16'b0000000000000000;
		15'h1738: char_row_bitmap <= 16'b0000000000000000;
		15'h1739: char_row_bitmap <= 16'b0000000000000000;
		15'h173a: char_row_bitmap <= 16'b0000000000000000;
		15'h173b: char_row_bitmap <= 16'b0000000000000000;
		15'h173c: char_row_bitmap <= 16'b0000000000000000;
		15'h173d: char_row_bitmap <= 16'b0000000000000000;
		15'h173e: char_row_bitmap <= 16'b0000000000000000;
		15'h173f: char_row_bitmap <= 16'b0000000000000000;
		15'h1740: char_row_bitmap <= 16'b0000000000000000;
		15'h1741: char_row_bitmap <= 16'b0000000000000000;
		15'h1742: char_row_bitmap <= 16'b0000000000000000;
		15'h1743: char_row_bitmap <= 16'b0000000000000000;
		15'h1744: char_row_bitmap <= 16'b0000000000000000;
		15'h1745: char_row_bitmap <= 16'b0000000000000000;
		15'h1746: char_row_bitmap <= 16'b0000000000000000;
		15'h1747: char_row_bitmap <= 16'b0000000000000000;
		15'h1748: char_row_bitmap <= 16'b0000000000000000;
		15'h1749: char_row_bitmap <= 16'b0000000000000000;
		15'h174a: char_row_bitmap <= 16'b0000000000000000;
		15'h174b: char_row_bitmap <= 16'b0000000000000000;
		15'h174c: char_row_bitmap <= 16'b0000000000000000;
		15'h174d: char_row_bitmap <= 16'b0000000000000000;
		15'h174e: char_row_bitmap <= 16'b0000000000000000;
		15'h174f: char_row_bitmap <= 16'b0000000000000000;
		15'h1750: char_row_bitmap <= 16'b0000000000000000;
		15'h1751: char_row_bitmap <= 16'b0000000000000000;
		15'h1752: char_row_bitmap <= 16'b0000000000000000;
		15'h1753: char_row_bitmap <= 16'b0000000000000000;
		15'h1754: char_row_bitmap <= 16'b0000000000000000;
		15'h1755: char_row_bitmap <= 16'b0000000000000000;
		15'h1756: char_row_bitmap <= 16'b0000000000000000;
		15'h1757: char_row_bitmap <= 16'b0000000000000000;
		15'h1758: char_row_bitmap <= 16'b0000000000000000;
		15'h1759: char_row_bitmap <= 16'b0000000000000000;
		15'h175a: char_row_bitmap <= 16'b0000000000000000;
		15'h175b: char_row_bitmap <= 16'b0000000000000000;
		15'h175c: char_row_bitmap <= 16'b0000000000000000;
		15'h175d: char_row_bitmap <= 16'b0000000000000000;
		15'h175e: char_row_bitmap <= 16'b0000000000000000;
		15'h175f: char_row_bitmap <= 16'b0000000000000000;
		15'h1760: char_row_bitmap <= 16'b0000000000000000;
		15'h1761: char_row_bitmap <= 16'b0000000000000000;
		15'h1762: char_row_bitmap <= 16'b0000000000000000;
		15'h1763: char_row_bitmap <= 16'b0000000000000000;
		15'h1764: char_row_bitmap <= 16'b0000000000000000;
		15'h1765: char_row_bitmap <= 16'b0000000000000000;
		15'h1766: char_row_bitmap <= 16'b0000000000000000;
		15'h1767: char_row_bitmap <= 16'b0000000000000000;
		15'h1768: char_row_bitmap <= 16'b0000000000000000;
		15'h1769: char_row_bitmap <= 16'b0000000000000000;
		15'h176a: char_row_bitmap <= 16'b0000000000000000;
		15'h176b: char_row_bitmap <= 16'b0000000000000000;
		15'h176c: char_row_bitmap <= 16'b0000000000000000;
		15'h176d: char_row_bitmap <= 16'b0000000000000000;
		15'h176e: char_row_bitmap <= 16'b0000000000000000;
		15'h176f: char_row_bitmap <= 16'b0000000000000000;
		15'h1770: char_row_bitmap <= 16'b0000000000000000;
		15'h1771: char_row_bitmap <= 16'b0000000000000000;
		15'h1772: char_row_bitmap <= 16'b0000000000000000;
		15'h1773: char_row_bitmap <= 16'b0000000000000000;
		15'h1774: char_row_bitmap <= 16'b0000000000000000;
		15'h1775: char_row_bitmap <= 16'b0000000000000000;
		15'h1776: char_row_bitmap <= 16'b0000000000000000;
		15'h1777: char_row_bitmap <= 16'b0000000000000000;
		15'h1778: char_row_bitmap <= 16'b0000000000000000;
		15'h1779: char_row_bitmap <= 16'b0000000000000000;
		15'h177a: char_row_bitmap <= 16'b0000000000000000;
		15'h177b: char_row_bitmap <= 16'b0000000000000000;
		15'h177c: char_row_bitmap <= 16'b0000000000000000;
		15'h177d: char_row_bitmap <= 16'b0000000000000000;
		15'h177e: char_row_bitmap <= 16'b0000000000000000;
		15'h177f: char_row_bitmap <= 16'b0000000000000000;
		15'h1780: char_row_bitmap <= 16'b0000000000000000;
		15'h1781: char_row_bitmap <= 16'b0000000000000000;
		15'h1782: char_row_bitmap <= 16'b0000000000000000;
		15'h1783: char_row_bitmap <= 16'b0000000000000000;
		15'h1784: char_row_bitmap <= 16'b0000000000000000;
		15'h1785: char_row_bitmap <= 16'b0000000000000000;
		15'h1786: char_row_bitmap <= 16'b0000000000000000;
		15'h1787: char_row_bitmap <= 16'b0000000000000000;
		15'h1788: char_row_bitmap <= 16'b0000000000000000;
		15'h1789: char_row_bitmap <= 16'b0000000000000000;
		15'h178a: char_row_bitmap <= 16'b0000000000000000;
		15'h178b: char_row_bitmap <= 16'b0000000000000000;
		15'h178c: char_row_bitmap <= 16'b0000000000000000;
		15'h178d: char_row_bitmap <= 16'b0000000000000000;
		15'h178e: char_row_bitmap <= 16'b0000000000000000;
		15'h178f: char_row_bitmap <= 16'b0000000000000000;
		15'h1790: char_row_bitmap <= 16'b0000000000000000;
		15'h1791: char_row_bitmap <= 16'b0000000000000000;
		15'h1792: char_row_bitmap <= 16'b0000000000000000;
		15'h1793: char_row_bitmap <= 16'b0000000000000000;
		15'h1794: char_row_bitmap <= 16'b0000000000000000;
		15'h1795: char_row_bitmap <= 16'b0000000000000000;
		15'h1796: char_row_bitmap <= 16'b0000000000000000;
		15'h1797: char_row_bitmap <= 16'b0000000000000000;
		15'h1798: char_row_bitmap <= 16'b0000000000000000;
		15'h1799: char_row_bitmap <= 16'b0000000000000000;
		15'h179a: char_row_bitmap <= 16'b0000000000000000;
		15'h179b: char_row_bitmap <= 16'b0000000000000000;
		15'h179c: char_row_bitmap <= 16'b0000000000000000;
		15'h179d: char_row_bitmap <= 16'b0000000000000000;
		15'h179e: char_row_bitmap <= 16'b0000000000000000;
		15'h179f: char_row_bitmap <= 16'b0000000000000000;
		15'h17a0: char_row_bitmap <= 16'b0000000000000000;
		15'h17a1: char_row_bitmap <= 16'b0000000000000000;
		15'h17a2: char_row_bitmap <= 16'b0000000000000000;
		15'h17a3: char_row_bitmap <= 16'b0000000000000000;
		15'h17a4: char_row_bitmap <= 16'b0000000000000000;
		15'h17a5: char_row_bitmap <= 16'b0000000000000000;
		15'h17a6: char_row_bitmap <= 16'b0000000000000000;
		15'h17a7: char_row_bitmap <= 16'b0000000000000000;
		15'h17a8: char_row_bitmap <= 16'b0000000000000000;
		15'h17a9: char_row_bitmap <= 16'b0000000000000000;
		15'h17aa: char_row_bitmap <= 16'b0000000000000000;
		15'h17ab: char_row_bitmap <= 16'b0000000000000000;
		15'h17ac: char_row_bitmap <= 16'b0000000000000000;
		15'h17ad: char_row_bitmap <= 16'b0000000000000000;
		15'h17ae: char_row_bitmap <= 16'b0000000000000000;
		15'h17af: char_row_bitmap <= 16'b0000000000000000;
		15'h17b0: char_row_bitmap <= 16'b0000000000000000;
		15'h17b1: char_row_bitmap <= 16'b0000000000000000;
		15'h17b2: char_row_bitmap <= 16'b0000000000000000;
		15'h17b3: char_row_bitmap <= 16'b0000000000000000;
		15'h17b4: char_row_bitmap <= 16'b0000000000000000;
		15'h17b5: char_row_bitmap <= 16'b0000000000000000;
		15'h17b6: char_row_bitmap <= 16'b0000000000000000;
		15'h17b7: char_row_bitmap <= 16'b0000000000000000;
		15'h17b8: char_row_bitmap <= 16'b0000000000000000;
		15'h17b9: char_row_bitmap <= 16'b0000000000000000;
		15'h17ba: char_row_bitmap <= 16'b0000000000000000;
		15'h17bb: char_row_bitmap <= 16'b0000000000000000;
		15'h17bc: char_row_bitmap <= 16'b0000000000000000;
		15'h17bd: char_row_bitmap <= 16'b0000000000000000;
		15'h17be: char_row_bitmap <= 16'b0000000000000000;
		15'h17bf: char_row_bitmap <= 16'b0000000000000000;
		15'h17c0: char_row_bitmap <= 16'b0000000000000000;
		15'h17c1: char_row_bitmap <= 16'b0000000000000000;
		15'h17c2: char_row_bitmap <= 16'b0000000000000000;
		15'h17c3: char_row_bitmap <= 16'b0000000000000000;
		15'h17c4: char_row_bitmap <= 16'b0000000000000000;
		15'h17c5: char_row_bitmap <= 16'b0000000000000000;
		15'h17c6: char_row_bitmap <= 16'b0000000000000000;
		15'h17c7: char_row_bitmap <= 16'b0000000000000000;
		15'h17c8: char_row_bitmap <= 16'b0000000000000000;
		15'h17c9: char_row_bitmap <= 16'b0000000000000000;
		15'h17ca: char_row_bitmap <= 16'b0000000000000000;
		15'h17cb: char_row_bitmap <= 16'b0000000000000000;
		15'h17cc: char_row_bitmap <= 16'b0000000000000000;
		15'h17cd: char_row_bitmap <= 16'b0000000000000000;
		15'h17ce: char_row_bitmap <= 16'b0000000000000000;
		15'h17cf: char_row_bitmap <= 16'b0000000000000000;
		15'h17d0: char_row_bitmap <= 16'b0000000000000000;
		15'h17d1: char_row_bitmap <= 16'b0000000000000000;
		15'h17d2: char_row_bitmap <= 16'b0000000000000000;
		15'h17d3: char_row_bitmap <= 16'b0000000000000000;
		15'h17d4: char_row_bitmap <= 16'b0000000000000000;
		15'h17d5: char_row_bitmap <= 16'b0000000000000000;
		15'h17d6: char_row_bitmap <= 16'b0000000000000000;
		15'h17d7: char_row_bitmap <= 16'b0000000000000000;
		15'h17d8: char_row_bitmap <= 16'b0000000000000000;
		15'h17d9: char_row_bitmap <= 16'b0000000000000000;
		15'h17da: char_row_bitmap <= 16'b0000000000000000;
		15'h17db: char_row_bitmap <= 16'b0000000000000000;
		15'h17dc: char_row_bitmap <= 16'b0000000000000000;
		15'h17dd: char_row_bitmap <= 16'b0000000000000000;
		15'h17de: char_row_bitmap <= 16'b0000000000000000;
		15'h17df: char_row_bitmap <= 16'b0000000000000000;
		15'h17e0: char_row_bitmap <= 16'b0000000000000000;
		15'h17e1: char_row_bitmap <= 16'b0000000000000000;
		15'h17e2: char_row_bitmap <= 16'b0000000000000000;
		15'h17e3: char_row_bitmap <= 16'b0000000000000000;
		15'h17e4: char_row_bitmap <= 16'b0000000000000000;
		15'h17e5: char_row_bitmap <= 16'b0000000000000000;
		15'h17e6: char_row_bitmap <= 16'b0000000000000000;
		15'h17e7: char_row_bitmap <= 16'b0000000000000000;
		15'h17e8: char_row_bitmap <= 16'b0000000000000000;
		15'h17e9: char_row_bitmap <= 16'b0000000000000000;
		15'h17ea: char_row_bitmap <= 16'b0000000000000000;
		15'h17eb: char_row_bitmap <= 16'b0000000000000000;
		15'h17ec: char_row_bitmap <= 16'b0000000000000000;
		15'h17ed: char_row_bitmap <= 16'b0000000000000000;
		15'h17ee: char_row_bitmap <= 16'b0000000000000000;
		15'h17ef: char_row_bitmap <= 16'b0000000000000000;
		15'h17f0: char_row_bitmap <= 16'b0000000000000000;
		15'h17f1: char_row_bitmap <= 16'b0000000000000000;
		15'h17f2: char_row_bitmap <= 16'b0000000000000000;
		15'h17f3: char_row_bitmap <= 16'b0000000000000000;
		15'h17f4: char_row_bitmap <= 16'b0000000000000000;
		15'h17f5: char_row_bitmap <= 16'b0000000000000000;
		15'h17f6: char_row_bitmap <= 16'b0000000000000000;
		15'h17f7: char_row_bitmap <= 16'b0000000000000000;
		15'h17f8: char_row_bitmap <= 16'b0000000000000000;
		15'h17f9: char_row_bitmap <= 16'b0000000000000000;
		15'h17fa: char_row_bitmap <= 16'b0000000000000000;
		15'h17fb: char_row_bitmap <= 16'b0000000000000000;
		15'h17fc: char_row_bitmap <= 16'b0000000000000000;
		15'h17fd: char_row_bitmap <= 16'b0000000000000000;
		15'h17fe: char_row_bitmap <= 16'b0000000000000000;
		15'h17ff: char_row_bitmap <= 16'b0000000000000000;
		15'h1800: char_row_bitmap <= 16'b0000000000000000;
		15'h1801: char_row_bitmap <= 16'b0000000000000000;
		15'h1802: char_row_bitmap <= 16'b0000000000000000;
		15'h1803: char_row_bitmap <= 16'b0000000000000000;
		15'h1804: char_row_bitmap <= 16'b0000000000000000;
		15'h1805: char_row_bitmap <= 16'b0000000000000000;
		15'h1806: char_row_bitmap <= 16'b0000000000000000;
		15'h1807: char_row_bitmap <= 16'b0000000000000000;
		15'h1808: char_row_bitmap <= 16'b0000000000000000;
		15'h1809: char_row_bitmap <= 16'b0000000000000000;
		15'h180a: char_row_bitmap <= 16'b0000000000000000;
		15'h180b: char_row_bitmap <= 16'b0000000000000000;
		15'h180c: char_row_bitmap <= 16'b0000000000000000;
		15'h180d: char_row_bitmap <= 16'b0000000000000000;
		15'h180e: char_row_bitmap <= 16'b0000000000000000;
		15'h180f: char_row_bitmap <= 16'b0000000000000000;
		15'h1810: char_row_bitmap <= 16'b0000000000000000;
		15'h1811: char_row_bitmap <= 16'b0000000000000000;
		15'h1812: char_row_bitmap <= 16'b0000000000000000;
		15'h1813: char_row_bitmap <= 16'b0000000000000000;
		15'h1814: char_row_bitmap <= 16'b0000000000000000;
		15'h1815: char_row_bitmap <= 16'b0000000000000000;
		15'h1816: char_row_bitmap <= 16'b0000000000000000;
		15'h1817: char_row_bitmap <= 16'b0000000000000000;
		15'h1818: char_row_bitmap <= 16'b0000000000000000;
		15'h1819: char_row_bitmap <= 16'b0000000000000000;
		15'h181a: char_row_bitmap <= 16'b0000000000000000;
		15'h181b: char_row_bitmap <= 16'b0000000000000000;
		15'h181c: char_row_bitmap <= 16'b0000000000000000;
		15'h181d: char_row_bitmap <= 16'b0000000000000000;
		15'h181e: char_row_bitmap <= 16'b0000000000000000;
		15'h181f: char_row_bitmap <= 16'b0000000000000000;
		15'h1820: char_row_bitmap <= 16'b0000000000000000;
		15'h1821: char_row_bitmap <= 16'b0000000000000000;
		15'h1822: char_row_bitmap <= 16'b0000000000000000;
		15'h1823: char_row_bitmap <= 16'b0000000000000000;
		15'h1824: char_row_bitmap <= 16'b0000000000000000;
		15'h1825: char_row_bitmap <= 16'b0000000000000000;
		15'h1826: char_row_bitmap <= 16'b0000000000000000;
		15'h1827: char_row_bitmap <= 16'b0000000000000000;
		15'h1828: char_row_bitmap <= 16'b0000000000000000;
		15'h1829: char_row_bitmap <= 16'b0000000000000000;
		15'h182a: char_row_bitmap <= 16'b0000000000000000;
		15'h182b: char_row_bitmap <= 16'b0000000000000000;
		15'h182c: char_row_bitmap <= 16'b0000000000000000;
		15'h182d: char_row_bitmap <= 16'b0000000000000000;
		15'h182e: char_row_bitmap <= 16'b0000000000000000;
		15'h182f: char_row_bitmap <= 16'b0000000000000000;
		15'h1830: char_row_bitmap <= 16'b0000000000000000;
		15'h1831: char_row_bitmap <= 16'b0000000000000000;
		15'h1832: char_row_bitmap <= 16'b0000000000000000;
		15'h1833: char_row_bitmap <= 16'b0000000000000000;
		15'h1834: char_row_bitmap <= 16'b0000000000000000;
		15'h1835: char_row_bitmap <= 16'b0000000000000000;
		15'h1836: char_row_bitmap <= 16'b0000000000000000;
		15'h1837: char_row_bitmap <= 16'b0000000000000000;
		15'h1838: char_row_bitmap <= 16'b0000000000000000;
		15'h1839: char_row_bitmap <= 16'b0000000000000000;
		15'h183a: char_row_bitmap <= 16'b0000000000000000;
		15'h183b: char_row_bitmap <= 16'b0000000000000000;
		15'h183c: char_row_bitmap <= 16'b0000000000000000;
		15'h183d: char_row_bitmap <= 16'b0000000000000000;
		15'h183e: char_row_bitmap <= 16'b0000000000000000;
		15'h183f: char_row_bitmap <= 16'b0000000000000000;
		15'h1840: char_row_bitmap <= 16'b0000000000000000;
		15'h1841: char_row_bitmap <= 16'b0000000000000000;
		15'h1842: char_row_bitmap <= 16'b0000000000000000;
		15'h1843: char_row_bitmap <= 16'b0000000000000000;
		15'h1844: char_row_bitmap <= 16'b0000000000000000;
		15'h1845: char_row_bitmap <= 16'b0000000000000000;
		15'h1846: char_row_bitmap <= 16'b0000000000000000;
		15'h1847: char_row_bitmap <= 16'b0000000000000000;
		15'h1848: char_row_bitmap <= 16'b0000000000000000;
		15'h1849: char_row_bitmap <= 16'b0000000000000000;
		15'h184a: char_row_bitmap <= 16'b0000000000000000;
		15'h184b: char_row_bitmap <= 16'b0000000000000000;
		15'h184c: char_row_bitmap <= 16'b0000000000000000;
		15'h184d: char_row_bitmap <= 16'b0000000000000000;
		15'h184e: char_row_bitmap <= 16'b0000000000000000;
		15'h184f: char_row_bitmap <= 16'b0000000000000000;
		15'h1850: char_row_bitmap <= 16'b0000000000000000;
		15'h1851: char_row_bitmap <= 16'b0000000000000000;
		15'h1852: char_row_bitmap <= 16'b0000000000000000;
		15'h1853: char_row_bitmap <= 16'b0000000000000000;
		15'h1854: char_row_bitmap <= 16'b0000000000000000;
		15'h1855: char_row_bitmap <= 16'b0000000000000000;
		15'h1856: char_row_bitmap <= 16'b0000000000000000;
		15'h1857: char_row_bitmap <= 16'b0000000000000000;
		15'h1858: char_row_bitmap <= 16'b0000000000000000;
		15'h1859: char_row_bitmap <= 16'b0000000000000000;
		15'h185a: char_row_bitmap <= 16'b0000000000000000;
		15'h185b: char_row_bitmap <= 16'b0000000000000000;
		15'h185c: char_row_bitmap <= 16'b0000000000000000;
		15'h185d: char_row_bitmap <= 16'b0000000000000000;
		15'h185e: char_row_bitmap <= 16'b0000000000000000;
		15'h185f: char_row_bitmap <= 16'b0000000000000000;
		15'h1860: char_row_bitmap <= 16'b0000000000000000;
		15'h1861: char_row_bitmap <= 16'b0000000000000000;
		15'h1862: char_row_bitmap <= 16'b0000000000000000;
		15'h1863: char_row_bitmap <= 16'b0000000000000000;
		15'h1864: char_row_bitmap <= 16'b0000000000000000;
		15'h1865: char_row_bitmap <= 16'b0000000000000000;
		15'h1866: char_row_bitmap <= 16'b0000000000000000;
		15'h1867: char_row_bitmap <= 16'b0000000000000000;
		15'h1868: char_row_bitmap <= 16'b0000000000000000;
		15'h1869: char_row_bitmap <= 16'b0000000000000000;
		15'h186a: char_row_bitmap <= 16'b0000000000000000;
		15'h186b: char_row_bitmap <= 16'b0000000000000000;
		15'h186c: char_row_bitmap <= 16'b0000000000000000;
		15'h186d: char_row_bitmap <= 16'b0000000000000000;
		15'h186e: char_row_bitmap <= 16'b0000000000000000;
		15'h186f: char_row_bitmap <= 16'b0000000000000000;
		15'h1870: char_row_bitmap <= 16'b0000000000000000;
		15'h1871: char_row_bitmap <= 16'b0000000000000000;
		15'h1872: char_row_bitmap <= 16'b0000000000000000;
		15'h1873: char_row_bitmap <= 16'b0000000000000000;
		15'h1874: char_row_bitmap <= 16'b0000000000000000;
		15'h1875: char_row_bitmap <= 16'b0000000000000000;
		15'h1876: char_row_bitmap <= 16'b0000000000000000;
		15'h1877: char_row_bitmap <= 16'b0000000000000000;
		15'h1878: char_row_bitmap <= 16'b0000000000000000;
		15'h1879: char_row_bitmap <= 16'b0000000000000000;
		15'h187a: char_row_bitmap <= 16'b0000000000000000;
		15'h187b: char_row_bitmap <= 16'b0000000000000000;
		15'h187c: char_row_bitmap <= 16'b0000000000000000;
		15'h187d: char_row_bitmap <= 16'b0000000000000000;
		15'h187e: char_row_bitmap <= 16'b0000000000000000;
		15'h187f: char_row_bitmap <= 16'b0000000000000000;
		15'h1880: char_row_bitmap <= 16'b0000000000000000;
		15'h1881: char_row_bitmap <= 16'b0000000000000000;
		15'h1882: char_row_bitmap <= 16'b0000000000000000;
		15'h1883: char_row_bitmap <= 16'b0000000000000000;
		15'h1884: char_row_bitmap <= 16'b0000000000000000;
		15'h1885: char_row_bitmap <= 16'b0000000000000000;
		15'h1886: char_row_bitmap <= 16'b0000000000000000;
		15'h1887: char_row_bitmap <= 16'b0000000000000000;
		15'h1888: char_row_bitmap <= 16'b0000000000000000;
		15'h1889: char_row_bitmap <= 16'b0000000000000000;
		15'h188a: char_row_bitmap <= 16'b0000000000000000;
		15'h188b: char_row_bitmap <= 16'b0000000000000000;
		15'h188c: char_row_bitmap <= 16'b0000000000000000;
		15'h188d: char_row_bitmap <= 16'b0000000000000000;
		15'h188e: char_row_bitmap <= 16'b0000000000000000;
		15'h188f: char_row_bitmap <= 16'b0000000000000000;
		15'h1890: char_row_bitmap <= 16'b0000000000000000;
		15'h1891: char_row_bitmap <= 16'b0000000000000000;
		15'h1892: char_row_bitmap <= 16'b0000000000000000;
		15'h1893: char_row_bitmap <= 16'b0000000000000000;
		15'h1894: char_row_bitmap <= 16'b0000000000000000;
		15'h1895: char_row_bitmap <= 16'b0000000000000000;
		15'h1896: char_row_bitmap <= 16'b0000000000000000;
		15'h1897: char_row_bitmap <= 16'b0000000000000000;
		15'h1898: char_row_bitmap <= 16'b0000000000000000;
		15'h1899: char_row_bitmap <= 16'b0000000000000000;
		15'h189a: char_row_bitmap <= 16'b0000000000000000;
		15'h189b: char_row_bitmap <= 16'b0000000000000000;
		15'h189c: char_row_bitmap <= 16'b0000000000000000;
		15'h189d: char_row_bitmap <= 16'b0000000000000000;
		15'h189e: char_row_bitmap <= 16'b0000000000000000;
		15'h189f: char_row_bitmap <= 16'b0000000000000000;
		15'h18a0: char_row_bitmap <= 16'b0000000000000000;
		15'h18a1: char_row_bitmap <= 16'b0000000000000000;
		15'h18a2: char_row_bitmap <= 16'b0000000000000000;
		15'h18a3: char_row_bitmap <= 16'b0000000000000000;
		15'h18a4: char_row_bitmap <= 16'b0000000000000000;
		15'h18a5: char_row_bitmap <= 16'b0000000000000000;
		15'h18a6: char_row_bitmap <= 16'b0000000000000000;
		15'h18a7: char_row_bitmap <= 16'b0000000000000000;
		15'h18a8: char_row_bitmap <= 16'b0000000000000000;
		15'h18a9: char_row_bitmap <= 16'b0000000000000000;
		15'h18aa: char_row_bitmap <= 16'b0000000000000000;
		15'h18ab: char_row_bitmap <= 16'b0000000000000000;
		15'h18ac: char_row_bitmap <= 16'b0000000000000000;
		15'h18ad: char_row_bitmap <= 16'b0000000000000000;
		15'h18ae: char_row_bitmap <= 16'b0000000000000000;
		15'h18af: char_row_bitmap <= 16'b0000000000000000;
		15'h18b0: char_row_bitmap <= 16'b0000000000000000;
		15'h18b1: char_row_bitmap <= 16'b0000000000000000;
		15'h18b2: char_row_bitmap <= 16'b0000000000000000;
		15'h18b3: char_row_bitmap <= 16'b0000000000000000;
		15'h18b4: char_row_bitmap <= 16'b0000000000000000;
		15'h18b5: char_row_bitmap <= 16'b0000000000000000;
		15'h18b6: char_row_bitmap <= 16'b0000000000000000;
		15'h18b7: char_row_bitmap <= 16'b0000000000000000;
		15'h18b8: char_row_bitmap <= 16'b0000000000000000;
		15'h18b9: char_row_bitmap <= 16'b0000000000000000;
		15'h18ba: char_row_bitmap <= 16'b0000000000000000;
		15'h18bb: char_row_bitmap <= 16'b0000000000000000;
		15'h18bc: char_row_bitmap <= 16'b0000000000000000;
		15'h18bd: char_row_bitmap <= 16'b0000000000000000;
		15'h18be: char_row_bitmap <= 16'b0000000000000000;
		15'h18bf: char_row_bitmap <= 16'b0000000000000000;
		15'h18c0: char_row_bitmap <= 16'b0000000000000000;
		15'h18c1: char_row_bitmap <= 16'b0000000000000000;
		15'h18c2: char_row_bitmap <= 16'b0000000000000000;
		15'h18c3: char_row_bitmap <= 16'b0000000000000000;
		15'h18c4: char_row_bitmap <= 16'b0000000000000000;
		15'h18c5: char_row_bitmap <= 16'b0000000000000000;
		15'h18c6: char_row_bitmap <= 16'b0000000000000000;
		15'h18c7: char_row_bitmap <= 16'b0000000000000000;
		15'h18c8: char_row_bitmap <= 16'b0000000000000000;
		15'h18c9: char_row_bitmap <= 16'b0000000000000000;
		15'h18ca: char_row_bitmap <= 16'b0000000000000000;
		15'h18cb: char_row_bitmap <= 16'b0000000000000000;
		15'h18cc: char_row_bitmap <= 16'b0000000000000000;
		15'h18cd: char_row_bitmap <= 16'b0000000000000000;
		15'h18ce: char_row_bitmap <= 16'b0000000000000000;
		15'h18cf: char_row_bitmap <= 16'b0000000000000000;
		15'h18d0: char_row_bitmap <= 16'b0000000000000000;
		15'h18d1: char_row_bitmap <= 16'b0000000000000000;
		15'h18d2: char_row_bitmap <= 16'b0000000000000000;
		15'h18d3: char_row_bitmap <= 16'b0000000000000000;
		15'h18d4: char_row_bitmap <= 16'b0000000000000000;
		15'h18d5: char_row_bitmap <= 16'b0000000000000000;
		15'h18d6: char_row_bitmap <= 16'b0000000000000000;
		15'h18d7: char_row_bitmap <= 16'b0000000000000000;
		15'h18d8: char_row_bitmap <= 16'b0000000000000000;
		15'h18d9: char_row_bitmap <= 16'b0000000000000000;
		15'h18da: char_row_bitmap <= 16'b0000000000000000;
		15'h18db: char_row_bitmap <= 16'b0000000000000000;
		15'h18dc: char_row_bitmap <= 16'b0000000000000000;
		15'h18dd: char_row_bitmap <= 16'b0000000000000000;
		15'h18de: char_row_bitmap <= 16'b0000000000000000;
		15'h18df: char_row_bitmap <= 16'b0000000000000000;
		15'h18e0: char_row_bitmap <= 16'b0000000000000000;
		15'h18e1: char_row_bitmap <= 16'b0000000000000000;
		15'h18e2: char_row_bitmap <= 16'b0000000000000000;
		15'h18e3: char_row_bitmap <= 16'b0000000000000000;
		15'h18e4: char_row_bitmap <= 16'b0000000000000000;
		15'h18e5: char_row_bitmap <= 16'b0000000000000000;
		15'h18e6: char_row_bitmap <= 16'b0000000000000000;
		15'h18e7: char_row_bitmap <= 16'b0000000000000000;
		15'h18e8: char_row_bitmap <= 16'b0000000000000000;
		15'h18e9: char_row_bitmap <= 16'b0000000000000000;
		15'h18ea: char_row_bitmap <= 16'b0000000000000000;
		15'h18eb: char_row_bitmap <= 16'b0000000000000000;
		15'h18ec: char_row_bitmap <= 16'b0000000000000000;
		15'h18ed: char_row_bitmap <= 16'b0000000000000000;
		15'h18ee: char_row_bitmap <= 16'b0000000000000000;
		15'h18ef: char_row_bitmap <= 16'b0000000000000000;
		15'h18f0: char_row_bitmap <= 16'b0000000000000000;
		15'h18f1: char_row_bitmap <= 16'b0000000000000000;
		15'h18f2: char_row_bitmap <= 16'b0000000000000000;
		15'h18f3: char_row_bitmap <= 16'b0000000000000000;
		15'h18f4: char_row_bitmap <= 16'b0000000000000000;
		15'h18f5: char_row_bitmap <= 16'b0000000000000000;
		15'h18f6: char_row_bitmap <= 16'b0000000000000000;
		15'h18f7: char_row_bitmap <= 16'b0000000000000000;
		15'h18f8: char_row_bitmap <= 16'b0000000000000000;
		15'h18f9: char_row_bitmap <= 16'b0000000000000000;
		15'h18fa: char_row_bitmap <= 16'b0000000000000000;
		15'h18fb: char_row_bitmap <= 16'b0000000000000000;
		15'h18fc: char_row_bitmap <= 16'b0000000000000000;
		15'h18fd: char_row_bitmap <= 16'b0000000000000000;
		15'h18fe: char_row_bitmap <= 16'b0000000000000000;
		15'h18ff: char_row_bitmap <= 16'b0000000000000000;
		15'h1900: char_row_bitmap <= 16'b0000000000000000;
		15'h1901: char_row_bitmap <= 16'b0000000000000000;
		15'h1902: char_row_bitmap <= 16'b0000000000000000;
		15'h1903: char_row_bitmap <= 16'b0000000000000000;
		15'h1904: char_row_bitmap <= 16'b0000000000000000;
		15'h1905: char_row_bitmap <= 16'b0000000000000000;
		15'h1906: char_row_bitmap <= 16'b0000000000000000;
		15'h1907: char_row_bitmap <= 16'b0000000000000000;
		15'h1908: char_row_bitmap <= 16'b0000000000000000;
		15'h1909: char_row_bitmap <= 16'b0000000000000000;
		15'h190a: char_row_bitmap <= 16'b0000000000000000;
		15'h190b: char_row_bitmap <= 16'b0000000000000000;
		15'h190c: char_row_bitmap <= 16'b0000000000000000;
		15'h190d: char_row_bitmap <= 16'b0000000000000000;
		15'h190e: char_row_bitmap <= 16'b0000000000000000;
		15'h190f: char_row_bitmap <= 16'b0000000000000000;
		15'h1910: char_row_bitmap <= 16'b0000000000000000;
		15'h1911: char_row_bitmap <= 16'b0000000000000000;
		15'h1912: char_row_bitmap <= 16'b0000000000000000;
		15'h1913: char_row_bitmap <= 16'b0000000000000000;
		15'h1914: char_row_bitmap <= 16'b0000000000000000;
		15'h1915: char_row_bitmap <= 16'b0000000000000000;
		15'h1916: char_row_bitmap <= 16'b0000000000000000;
		15'h1917: char_row_bitmap <= 16'b0000000000000000;
		15'h1918: char_row_bitmap <= 16'b0000000000000000;
		15'h1919: char_row_bitmap <= 16'b0000000000000000;
		15'h191a: char_row_bitmap <= 16'b0000000000000000;
		15'h191b: char_row_bitmap <= 16'b0000000000000000;
		15'h191c: char_row_bitmap <= 16'b0000000000000000;
		15'h191d: char_row_bitmap <= 16'b0000000000000000;
		15'h191e: char_row_bitmap <= 16'b0000000000000000;
		15'h191f: char_row_bitmap <= 16'b0000000000000000;
		15'h1920: char_row_bitmap <= 16'b0000000000000000;
		15'h1921: char_row_bitmap <= 16'b0000000000000000;
		15'h1922: char_row_bitmap <= 16'b0000000000000000;
		15'h1923: char_row_bitmap <= 16'b0000000000000000;
		15'h1924: char_row_bitmap <= 16'b0000000000000000;
		15'h1925: char_row_bitmap <= 16'b0000000000000000;
		15'h1926: char_row_bitmap <= 16'b0000000000000000;
		15'h1927: char_row_bitmap <= 16'b0000000000000000;
		15'h1928: char_row_bitmap <= 16'b0000000000000000;
		15'h1929: char_row_bitmap <= 16'b0000000000000000;
		15'h192a: char_row_bitmap <= 16'b0000000000000000;
		15'h192b: char_row_bitmap <= 16'b0000000000000000;
		15'h192c: char_row_bitmap <= 16'b0000000000000000;
		15'h192d: char_row_bitmap <= 16'b0000000000000000;
		15'h192e: char_row_bitmap <= 16'b0000000000000000;
		15'h192f: char_row_bitmap <= 16'b0000000000000000;
		15'h1930: char_row_bitmap <= 16'b0000000000000000;
		15'h1931: char_row_bitmap <= 16'b0000000000000000;
		15'h1932: char_row_bitmap <= 16'b0000000000000000;
		15'h1933: char_row_bitmap <= 16'b0000000000000000;
		15'h1934: char_row_bitmap <= 16'b0000000000000000;
		15'h1935: char_row_bitmap <= 16'b0000000000000000;
		15'h1936: char_row_bitmap <= 16'b0000000000000000;
		15'h1937: char_row_bitmap <= 16'b0000000000000000;
		15'h1938: char_row_bitmap <= 16'b0000000000000000;
		15'h1939: char_row_bitmap <= 16'b0000000000000000;
		15'h193a: char_row_bitmap <= 16'b0000000000000000;
		15'h193b: char_row_bitmap <= 16'b0000000000000000;
		15'h193c: char_row_bitmap <= 16'b0000000000000000;
		15'h193d: char_row_bitmap <= 16'b0000000000000000;
		15'h193e: char_row_bitmap <= 16'b0000000000000000;
		15'h193f: char_row_bitmap <= 16'b0000000000000000;
		15'h1940: char_row_bitmap <= 16'b0000000000000000;
		15'h1941: char_row_bitmap <= 16'b0000000000000000;
		15'h1942: char_row_bitmap <= 16'b0000000000000000;
		15'h1943: char_row_bitmap <= 16'b0000000000000000;
		15'h1944: char_row_bitmap <= 16'b0000000000000000;
		15'h1945: char_row_bitmap <= 16'b0000000000000000;
		15'h1946: char_row_bitmap <= 16'b0000000000000000;
		15'h1947: char_row_bitmap <= 16'b0000000000000000;
		15'h1948: char_row_bitmap <= 16'b0000000000000000;
		15'h1949: char_row_bitmap <= 16'b0000000000000000;
		15'h194a: char_row_bitmap <= 16'b0000000000000000;
		15'h194b: char_row_bitmap <= 16'b0000000000000000;
		15'h194c: char_row_bitmap <= 16'b0000000000000000;
		15'h194d: char_row_bitmap <= 16'b0000000000000000;
		15'h194e: char_row_bitmap <= 16'b0000000000000000;
		15'h194f: char_row_bitmap <= 16'b0000000000000000;
		15'h1950: char_row_bitmap <= 16'b0000000000000000;
		15'h1951: char_row_bitmap <= 16'b0000000000000000;
		15'h1952: char_row_bitmap <= 16'b0000000000000000;
		15'h1953: char_row_bitmap <= 16'b0000000000000000;
		15'h1954: char_row_bitmap <= 16'b0000000000000000;
		15'h1955: char_row_bitmap <= 16'b0000000000000000;
		15'h1956: char_row_bitmap <= 16'b0000000000000000;
		15'h1957: char_row_bitmap <= 16'b0000000000000000;
		15'h1958: char_row_bitmap <= 16'b0000000000000000;
		15'h1959: char_row_bitmap <= 16'b0000000000000000;
		15'h195a: char_row_bitmap <= 16'b0000000000000000;
		15'h195b: char_row_bitmap <= 16'b0000000000000000;
		15'h195c: char_row_bitmap <= 16'b0000000000000000;
		15'h195d: char_row_bitmap <= 16'b0000000000000000;
		15'h195e: char_row_bitmap <= 16'b0000000000000000;
		15'h195f: char_row_bitmap <= 16'b0000000000000000;
		15'h1960: char_row_bitmap <= 16'b0000000000000000;
		15'h1961: char_row_bitmap <= 16'b0000000000000000;
		15'h1962: char_row_bitmap <= 16'b0000000000000000;
		15'h1963: char_row_bitmap <= 16'b0000000000000000;
		15'h1964: char_row_bitmap <= 16'b0000000000000000;
		15'h1965: char_row_bitmap <= 16'b0000000000000000;
		15'h1966: char_row_bitmap <= 16'b0000000000000000;
		15'h1967: char_row_bitmap <= 16'b0000000000000000;
		15'h1968: char_row_bitmap <= 16'b0000000000000000;
		15'h1969: char_row_bitmap <= 16'b0000000000000000;
		15'h196a: char_row_bitmap <= 16'b0000000000000000;
		15'h196b: char_row_bitmap <= 16'b0000000000000000;
		15'h196c: char_row_bitmap <= 16'b0000000000000000;
		15'h196d: char_row_bitmap <= 16'b0000000000000000;
		15'h196e: char_row_bitmap <= 16'b0000000000000000;
		15'h196f: char_row_bitmap <= 16'b0000000000000000;
		15'h1970: char_row_bitmap <= 16'b0000000000000000;
		15'h1971: char_row_bitmap <= 16'b0000000000000000;
		15'h1972: char_row_bitmap <= 16'b0000000000000000;
		15'h1973: char_row_bitmap <= 16'b0000000000000000;
		15'h1974: char_row_bitmap <= 16'b0000000000000000;
		15'h1975: char_row_bitmap <= 16'b0000000000000000;
		15'h1976: char_row_bitmap <= 16'b0000000000000000;
		15'h1977: char_row_bitmap <= 16'b0000000000000000;
		15'h1978: char_row_bitmap <= 16'b0000000000000000;
		15'h1979: char_row_bitmap <= 16'b0000000000000000;
		15'h197a: char_row_bitmap <= 16'b0000000000000000;
		15'h197b: char_row_bitmap <= 16'b0000000000000000;
		15'h197c: char_row_bitmap <= 16'b0000000000000000;
		15'h197d: char_row_bitmap <= 16'b0000000000000000;
		15'h197e: char_row_bitmap <= 16'b0000000000000000;
		15'h197f: char_row_bitmap <= 16'b0000000000000000;
		15'h1980: char_row_bitmap <= 16'b0000000000000000;
		15'h1981: char_row_bitmap <= 16'b0000000000000000;
		15'h1982: char_row_bitmap <= 16'b0000000000000000;
		15'h1983: char_row_bitmap <= 16'b0000000000000000;
		15'h1984: char_row_bitmap <= 16'b0000000000000000;
		15'h1985: char_row_bitmap <= 16'b0000000000000000;
		15'h1986: char_row_bitmap <= 16'b0000000000000000;
		15'h1987: char_row_bitmap <= 16'b0000000000000000;
		15'h1988: char_row_bitmap <= 16'b0000000000000000;
		15'h1989: char_row_bitmap <= 16'b0000000000000000;
		15'h198a: char_row_bitmap <= 16'b0000000000000000;
		15'h198b: char_row_bitmap <= 16'b0000000000000000;
		15'h198c: char_row_bitmap <= 16'b0000000000000000;
		15'h198d: char_row_bitmap <= 16'b0000000000000000;
		15'h198e: char_row_bitmap <= 16'b0000000000000000;
		15'h198f: char_row_bitmap <= 16'b0000000000000000;
		15'h1990: char_row_bitmap <= 16'b0000000000000000;
		15'h1991: char_row_bitmap <= 16'b0000000000000000;
		15'h1992: char_row_bitmap <= 16'b0000000000000000;
		15'h1993: char_row_bitmap <= 16'b0000000000000000;
		15'h1994: char_row_bitmap <= 16'b0000000000000000;
		15'h1995: char_row_bitmap <= 16'b0000000000000000;
		15'h1996: char_row_bitmap <= 16'b0000000000000000;
		15'h1997: char_row_bitmap <= 16'b0000000000000000;
		15'h1998: char_row_bitmap <= 16'b0000000000000000;
		15'h1999: char_row_bitmap <= 16'b0000000000000000;
		15'h199a: char_row_bitmap <= 16'b0000000000000000;
		15'h199b: char_row_bitmap <= 16'b0000000000000000;
		15'h199c: char_row_bitmap <= 16'b0000000000000000;
		15'h199d: char_row_bitmap <= 16'b0000000000000000;
		15'h199e: char_row_bitmap <= 16'b0000000000000000;
		15'h199f: char_row_bitmap <= 16'b0000000000000000;
		15'h19a0: char_row_bitmap <= 16'b0000000000000000;
		15'h19a1: char_row_bitmap <= 16'b0000000000000000;
		15'h19a2: char_row_bitmap <= 16'b0000000000000000;
		15'h19a3: char_row_bitmap <= 16'b0000000000000000;
		15'h19a4: char_row_bitmap <= 16'b0000000000000000;
		15'h19a5: char_row_bitmap <= 16'b0000000000000000;
		15'h19a6: char_row_bitmap <= 16'b0000000000000000;
		15'h19a7: char_row_bitmap <= 16'b0000000000000000;
		15'h19a8: char_row_bitmap <= 16'b0000000000000000;
		15'h19a9: char_row_bitmap <= 16'b0000000000000000;
		15'h19aa: char_row_bitmap <= 16'b0000000000000000;
		15'h19ab: char_row_bitmap <= 16'b0000000000000000;
		15'h19ac: char_row_bitmap <= 16'b0000000000000000;
		15'h19ad: char_row_bitmap <= 16'b0000000000000000;
		15'h19ae: char_row_bitmap <= 16'b0000000000000000;
		15'h19af: char_row_bitmap <= 16'b0000000000000000;
		15'h19b0: char_row_bitmap <= 16'b0000000000000000;
		15'h19b1: char_row_bitmap <= 16'b0000000000000000;
		15'h19b2: char_row_bitmap <= 16'b0000000000000000;
		15'h19b3: char_row_bitmap <= 16'b0000000000000000;
		15'h19b4: char_row_bitmap <= 16'b0000000000000000;
		15'h19b5: char_row_bitmap <= 16'b0000000000000000;
		15'h19b6: char_row_bitmap <= 16'b0000000000000000;
		15'h19b7: char_row_bitmap <= 16'b0000000000000000;
		15'h19b8: char_row_bitmap <= 16'b0000000000000000;
		15'h19b9: char_row_bitmap <= 16'b0000000000000000;
		15'h19ba: char_row_bitmap <= 16'b0000000000000000;
		15'h19bb: char_row_bitmap <= 16'b0000000000000000;
		15'h19bc: char_row_bitmap <= 16'b0000000000000000;
		15'h19bd: char_row_bitmap <= 16'b0000000000000000;
		15'h19be: char_row_bitmap <= 16'b0000000000000000;
		15'h19bf: char_row_bitmap <= 16'b0000000000000000;
		15'h19c0: char_row_bitmap <= 16'b0000000000000000;
		15'h19c1: char_row_bitmap <= 16'b0000000000000000;
		15'h19c2: char_row_bitmap <= 16'b0000000000000000;
		15'h19c3: char_row_bitmap <= 16'b0000000000000000;
		15'h19c4: char_row_bitmap <= 16'b0000000000000000;
		15'h19c5: char_row_bitmap <= 16'b0000000000000000;
		15'h19c6: char_row_bitmap <= 16'b0000000000000000;
		15'h19c7: char_row_bitmap <= 16'b0000000000000000;
		15'h19c8: char_row_bitmap <= 16'b0000000000000000;
		15'h19c9: char_row_bitmap <= 16'b0000000000000000;
		15'h19ca: char_row_bitmap <= 16'b0000000000000000;
		15'h19cb: char_row_bitmap <= 16'b0000000000000000;
		15'h19cc: char_row_bitmap <= 16'b0000000000000000;
		15'h19cd: char_row_bitmap <= 16'b0000000000000000;
		15'h19ce: char_row_bitmap <= 16'b0000000000000000;
		15'h19cf: char_row_bitmap <= 16'b0000000000000000;
		15'h19d0: char_row_bitmap <= 16'b0000000000000000;
		15'h19d1: char_row_bitmap <= 16'b0000000000000000;
		15'h19d2: char_row_bitmap <= 16'b0000000000000000;
		15'h19d3: char_row_bitmap <= 16'b0000000000000000;
		15'h19d4: char_row_bitmap <= 16'b0000000000000000;
		15'h19d5: char_row_bitmap <= 16'b0000000000000000;
		15'h19d6: char_row_bitmap <= 16'b0000000000000000;
		15'h19d7: char_row_bitmap <= 16'b0000000000000000;
		15'h19d8: char_row_bitmap <= 16'b0000000000000000;
		15'h19d9: char_row_bitmap <= 16'b0000000000000000;
		15'h19da: char_row_bitmap <= 16'b0000000000000000;
		15'h19db: char_row_bitmap <= 16'b0000000000000000;
		15'h19dc: char_row_bitmap <= 16'b0000000000000000;
		15'h19dd: char_row_bitmap <= 16'b0000000000000000;
		15'h19de: char_row_bitmap <= 16'b0000000000000000;
		15'h19df: char_row_bitmap <= 16'b0000000000000000;
		15'h19e0: char_row_bitmap <= 16'b0000000000000000;
		15'h19e1: char_row_bitmap <= 16'b0000000000000000;
		15'h19e2: char_row_bitmap <= 16'b0000000000000000;
		15'h19e3: char_row_bitmap <= 16'b0000000000000000;
		15'h19e4: char_row_bitmap <= 16'b0000000000000000;
		15'h19e5: char_row_bitmap <= 16'b0000000000000000;
		15'h19e6: char_row_bitmap <= 16'b0000000000000000;
		15'h19e7: char_row_bitmap <= 16'b0000000000000000;
		15'h19e8: char_row_bitmap <= 16'b0000000000000000;
		15'h19e9: char_row_bitmap <= 16'b0000000000000000;
		15'h19ea: char_row_bitmap <= 16'b0000000000000000;
		15'h19eb: char_row_bitmap <= 16'b0000000000000000;
		15'h19ec: char_row_bitmap <= 16'b0000000000000000;
		15'h19ed: char_row_bitmap <= 16'b0000000000000000;
		15'h19ee: char_row_bitmap <= 16'b0000000000000000;
		15'h19ef: char_row_bitmap <= 16'b0000000000000000;
		15'h19f0: char_row_bitmap <= 16'b0000000000000000;
		15'h19f1: char_row_bitmap <= 16'b0000000000000000;
		15'h19f2: char_row_bitmap <= 16'b0000000000000000;
		15'h19f3: char_row_bitmap <= 16'b0000000000000000;
		15'h19f4: char_row_bitmap <= 16'b0000000000000000;
		15'h19f5: char_row_bitmap <= 16'b0000000000000000;
		15'h19f6: char_row_bitmap <= 16'b0000000000000000;
		15'h19f7: char_row_bitmap <= 16'b0000000000000000;
		15'h19f8: char_row_bitmap <= 16'b0000000000000000;
		15'h19f9: char_row_bitmap <= 16'b0000000000000000;
		15'h19fa: char_row_bitmap <= 16'b0000000000000000;
		15'h19fb: char_row_bitmap <= 16'b0000000000000000;
		15'h19fc: char_row_bitmap <= 16'b0000000000000000;
		15'h19fd: char_row_bitmap <= 16'b0000000000000000;
		15'h19fe: char_row_bitmap <= 16'b0000000000000000;
		15'h19ff: char_row_bitmap <= 16'b0000000000000000;
		15'h1a00: char_row_bitmap <= 16'b0000000000000000;
		15'h1a01: char_row_bitmap <= 16'b0000000000000000;
		15'h1a02: char_row_bitmap <= 16'b0000000000000000;
		15'h1a03: char_row_bitmap <= 16'b0000000000000000;
		15'h1a04: char_row_bitmap <= 16'b0000000000000000;
		15'h1a05: char_row_bitmap <= 16'b0000000000000000;
		15'h1a06: char_row_bitmap <= 16'b0000000000000000;
		15'h1a07: char_row_bitmap <= 16'b0000000000000000;
		15'h1a08: char_row_bitmap <= 16'b0000000000000000;
		15'h1a09: char_row_bitmap <= 16'b0000000000000000;
		15'h1a0a: char_row_bitmap <= 16'b0000000000000000;
		15'h1a0b: char_row_bitmap <= 16'b0000000000000000;
		15'h1a0c: char_row_bitmap <= 16'b0000000000000000;
		15'h1a0d: char_row_bitmap <= 16'b0000000000000000;
		15'h1a0e: char_row_bitmap <= 16'b0000000000000000;
		15'h1a0f: char_row_bitmap <= 16'b0000000000000000;
		15'h1a10: char_row_bitmap <= 16'b0000000000000000;
		15'h1a11: char_row_bitmap <= 16'b0000000000000000;
		15'h1a12: char_row_bitmap <= 16'b0000000000000000;
		15'h1a13: char_row_bitmap <= 16'b0000000000000000;
		15'h1a14: char_row_bitmap <= 16'b0000000000000000;
		15'h1a15: char_row_bitmap <= 16'b0000000000000000;
		15'h1a16: char_row_bitmap <= 16'b0000000000000000;
		15'h1a17: char_row_bitmap <= 16'b0000000000000000;
		15'h1a18: char_row_bitmap <= 16'b0000000000000000;
		15'h1a19: char_row_bitmap <= 16'b0000000000000000;
		15'h1a1a: char_row_bitmap <= 16'b0000000000000000;
		15'h1a1b: char_row_bitmap <= 16'b0000000000000000;
		15'h1a1c: char_row_bitmap <= 16'b0000000000000000;
		15'h1a1d: char_row_bitmap <= 16'b0000000000000000;
		15'h1a1e: char_row_bitmap <= 16'b0000000000000000;
		15'h1a1f: char_row_bitmap <= 16'b0000000000000000;
		15'h1a20: char_row_bitmap <= 16'b0000000000000000;
		15'h1a21: char_row_bitmap <= 16'b0000000000000000;
		15'h1a22: char_row_bitmap <= 16'b0000000000000000;
		15'h1a23: char_row_bitmap <= 16'b0000000000000000;
		15'h1a24: char_row_bitmap <= 16'b0000000000000000;
		15'h1a25: char_row_bitmap <= 16'b0000000000000000;
		15'h1a26: char_row_bitmap <= 16'b0000000000000000;
		15'h1a27: char_row_bitmap <= 16'b0000000000000000;
		15'h1a28: char_row_bitmap <= 16'b0000000000000000;
		15'h1a29: char_row_bitmap <= 16'b0000000000000000;
		15'h1a2a: char_row_bitmap <= 16'b0000000000000000;
		15'h1a2b: char_row_bitmap <= 16'b0000000000000000;
		15'h1a2c: char_row_bitmap <= 16'b0000000000000000;
		15'h1a2d: char_row_bitmap <= 16'b0000000000000000;
		15'h1a2e: char_row_bitmap <= 16'b0000000000000000;
		15'h1a2f: char_row_bitmap <= 16'b0000000000000000;
		15'h1a30: char_row_bitmap <= 16'b0000000000000000;
		15'h1a31: char_row_bitmap <= 16'b0000000000000000;
		15'h1a32: char_row_bitmap <= 16'b0000000000000000;
		15'h1a33: char_row_bitmap <= 16'b0000000000000000;
		15'h1a34: char_row_bitmap <= 16'b0000000000000000;
		15'h1a35: char_row_bitmap <= 16'b0000000000000000;
		15'h1a36: char_row_bitmap <= 16'b0000000000000000;
		15'h1a37: char_row_bitmap <= 16'b0000000000000000;
		15'h1a38: char_row_bitmap <= 16'b0000000000000000;
		15'h1a39: char_row_bitmap <= 16'b0000000000000000;
		15'h1a3a: char_row_bitmap <= 16'b0000000000000000;
		15'h1a3b: char_row_bitmap <= 16'b0000000000000000;
		15'h1a3c: char_row_bitmap <= 16'b0000000000000000;
		15'h1a3d: char_row_bitmap <= 16'b0000000000000000;
		15'h1a3e: char_row_bitmap <= 16'b0000000000000000;
		15'h1a3f: char_row_bitmap <= 16'b0000000000000000;
		15'h1a40: char_row_bitmap <= 16'b0000000000000000;
		15'h1a41: char_row_bitmap <= 16'b0000000000000000;
		15'h1a42: char_row_bitmap <= 16'b0000000000000000;
		15'h1a43: char_row_bitmap <= 16'b0000000000000000;
		15'h1a44: char_row_bitmap <= 16'b0000000000000000;
		15'h1a45: char_row_bitmap <= 16'b0000000000000000;
		15'h1a46: char_row_bitmap <= 16'b0000000000000000;
		15'h1a47: char_row_bitmap <= 16'b0000000000000000;
		15'h1a48: char_row_bitmap <= 16'b0000000000000000;
		15'h1a49: char_row_bitmap <= 16'b0000000000000000;
		15'h1a4a: char_row_bitmap <= 16'b0000000000000000;
		15'h1a4b: char_row_bitmap <= 16'b0000000000000000;
		15'h1a4c: char_row_bitmap <= 16'b0000000000000000;
		15'h1a4d: char_row_bitmap <= 16'b0000000000000000;
		15'h1a4e: char_row_bitmap <= 16'b0000000000000000;
		15'h1a4f: char_row_bitmap <= 16'b0000000000000000;
		15'h1a50: char_row_bitmap <= 16'b0000000000000000;
		15'h1a51: char_row_bitmap <= 16'b0000000000000000;
		15'h1a52: char_row_bitmap <= 16'b0000000000000000;
		15'h1a53: char_row_bitmap <= 16'b0000000000000000;
		15'h1a54: char_row_bitmap <= 16'b0000000000000000;
		15'h1a55: char_row_bitmap <= 16'b0000000000000000;
		15'h1a56: char_row_bitmap <= 16'b0000000000000000;
		15'h1a57: char_row_bitmap <= 16'b0000000000000000;
		15'h1a58: char_row_bitmap <= 16'b0000000000000000;
		15'h1a59: char_row_bitmap <= 16'b0000000000000000;
		15'h1a5a: char_row_bitmap <= 16'b0000000000000000;
		15'h1a5b: char_row_bitmap <= 16'b0000000000000000;
		15'h1a5c: char_row_bitmap <= 16'b0000000000000000;
		15'h1a5d: char_row_bitmap <= 16'b0000000000000000;
		15'h1a5e: char_row_bitmap <= 16'b0000000000000000;
		15'h1a5f: char_row_bitmap <= 16'b0000000000000000;
		15'h1a60: char_row_bitmap <= 16'b0000000000000000;
		15'h1a61: char_row_bitmap <= 16'b0000000000000000;
		15'h1a62: char_row_bitmap <= 16'b0000000000000000;
		15'h1a63: char_row_bitmap <= 16'b0000000000000000;
		15'h1a64: char_row_bitmap <= 16'b0000000000000000;
		15'h1a65: char_row_bitmap <= 16'b0000000000000000;
		15'h1a66: char_row_bitmap <= 16'b0000000000000000;
		15'h1a67: char_row_bitmap <= 16'b0000000000000000;
		15'h1a68: char_row_bitmap <= 16'b0000000000000000;
		15'h1a69: char_row_bitmap <= 16'b0000000000000000;
		15'h1a6a: char_row_bitmap <= 16'b0000000000000000;
		15'h1a6b: char_row_bitmap <= 16'b0000000000000000;
		15'h1a6c: char_row_bitmap <= 16'b0000000000000000;
		15'h1a6d: char_row_bitmap <= 16'b0000000000000000;
		15'h1a6e: char_row_bitmap <= 16'b0000000000000000;
		15'h1a6f: char_row_bitmap <= 16'b0000000000000000;
		15'h1a70: char_row_bitmap <= 16'b0000000000000000;
		15'h1a71: char_row_bitmap <= 16'b0000000000000000;
		15'h1a72: char_row_bitmap <= 16'b0000000000000000;
		15'h1a73: char_row_bitmap <= 16'b0000000000000000;
		15'h1a74: char_row_bitmap <= 16'b0000000000000000;
		15'h1a75: char_row_bitmap <= 16'b0000000000000000;
		15'h1a76: char_row_bitmap <= 16'b0000000000000000;
		15'h1a77: char_row_bitmap <= 16'b0000000000000000;
		15'h1a78: char_row_bitmap <= 16'b0000000000000000;
		15'h1a79: char_row_bitmap <= 16'b0000000000000000;
		15'h1a7a: char_row_bitmap <= 16'b0000000000000000;
		15'h1a7b: char_row_bitmap <= 16'b0000000000000000;
		15'h1a7c: char_row_bitmap <= 16'b0000000000000000;
		15'h1a7d: char_row_bitmap <= 16'b0000000000000000;
		15'h1a7e: char_row_bitmap <= 16'b0000000000000000;
		15'h1a7f: char_row_bitmap <= 16'b0000000000000000;
		15'h1a80: char_row_bitmap <= 16'b0000000000000000;
		15'h1a81: char_row_bitmap <= 16'b0000000000000000;
		15'h1a82: char_row_bitmap <= 16'b0000000000000000;
		15'h1a83: char_row_bitmap <= 16'b0000000000000000;
		15'h1a84: char_row_bitmap <= 16'b0000000000000000;
		15'h1a85: char_row_bitmap <= 16'b0000000000000000;
		15'h1a86: char_row_bitmap <= 16'b0000000000000000;
		15'h1a87: char_row_bitmap <= 16'b0000000000000000;
		15'h1a88: char_row_bitmap <= 16'b0000000000000000;
		15'h1a89: char_row_bitmap <= 16'b0000000000000000;
		15'h1a8a: char_row_bitmap <= 16'b0000000000000000;
		15'h1a8b: char_row_bitmap <= 16'b0000000000000000;
		15'h1a8c: char_row_bitmap <= 16'b0000000000000000;
		15'h1a8d: char_row_bitmap <= 16'b0000000000000000;
		15'h1a8e: char_row_bitmap <= 16'b0000000000000000;
		15'h1a8f: char_row_bitmap <= 16'b0000000000000000;
		15'h1a90: char_row_bitmap <= 16'b0000000000000000;
		15'h1a91: char_row_bitmap <= 16'b0000000000000000;
		15'h1a92: char_row_bitmap <= 16'b0000000000000000;
		15'h1a93: char_row_bitmap <= 16'b0000000000000000;
		15'h1a94: char_row_bitmap <= 16'b0000000000000000;
		15'h1a95: char_row_bitmap <= 16'b0000000000000000;
		15'h1a96: char_row_bitmap <= 16'b0000000000000000;
		15'h1a97: char_row_bitmap <= 16'b0000000000000000;
		15'h1a98: char_row_bitmap <= 16'b0000000000000000;
		15'h1a99: char_row_bitmap <= 16'b0000000000000000;
		15'h1a9a: char_row_bitmap <= 16'b0000000000000000;
		15'h1a9b: char_row_bitmap <= 16'b0000000000000000;
		15'h1a9c: char_row_bitmap <= 16'b0000000000000000;
		15'h1a9d: char_row_bitmap <= 16'b0000000000000000;
		15'h1a9e: char_row_bitmap <= 16'b0000000000000000;
		15'h1a9f: char_row_bitmap <= 16'b0000000000000000;
		15'h1aa0: char_row_bitmap <= 16'b0000000000000000;
		15'h1aa1: char_row_bitmap <= 16'b0000000000000000;
		15'h1aa2: char_row_bitmap <= 16'b0000000000000000;
		15'h1aa3: char_row_bitmap <= 16'b0000000000000000;
		15'h1aa4: char_row_bitmap <= 16'b0000000000000000;
		15'h1aa5: char_row_bitmap <= 16'b0000000000000000;
		15'h1aa6: char_row_bitmap <= 16'b0000000000000000;
		15'h1aa7: char_row_bitmap <= 16'b0000000000000000;
		15'h1aa8: char_row_bitmap <= 16'b0000000000000000;
		15'h1aa9: char_row_bitmap <= 16'b0000000000000000;
		15'h1aaa: char_row_bitmap <= 16'b0000000000000000;
		15'h1aab: char_row_bitmap <= 16'b0000000000000000;
		15'h1aac: char_row_bitmap <= 16'b0000000000000000;
		15'h1aad: char_row_bitmap <= 16'b0000000000000000;
		15'h1aae: char_row_bitmap <= 16'b0000000000000000;
		15'h1aaf: char_row_bitmap <= 16'b0000000000000000;
		15'h1ab0: char_row_bitmap <= 16'b0000000000000000;
		15'h1ab1: char_row_bitmap <= 16'b0000000000000000;
		15'h1ab2: char_row_bitmap <= 16'b0000000000000000;
		15'h1ab3: char_row_bitmap <= 16'b0000000000000000;
		15'h1ab4: char_row_bitmap <= 16'b0000000000000000;
		15'h1ab5: char_row_bitmap <= 16'b0000000000000000;
		15'h1ab6: char_row_bitmap <= 16'b0000000000000000;
		15'h1ab7: char_row_bitmap <= 16'b0000000000000000;
		15'h1ab8: char_row_bitmap <= 16'b0000000000000000;
		15'h1ab9: char_row_bitmap <= 16'b0000000000000000;
		15'h1aba: char_row_bitmap <= 16'b0000000000000000;
		15'h1abb: char_row_bitmap <= 16'b0000000000000000;
		15'h1abc: char_row_bitmap <= 16'b0000000000000000;
		15'h1abd: char_row_bitmap <= 16'b0000000000000000;
		15'h1abe: char_row_bitmap <= 16'b0000000000000000;
		15'h1abf: char_row_bitmap <= 16'b0000000000000000;
		15'h1ac0: char_row_bitmap <= 16'b0000000000000000;
		15'h1ac1: char_row_bitmap <= 16'b0000000000000000;
		15'h1ac2: char_row_bitmap <= 16'b0000000000000000;
		15'h1ac3: char_row_bitmap <= 16'b0000000000000000;
		15'h1ac4: char_row_bitmap <= 16'b0000000000000000;
		15'h1ac5: char_row_bitmap <= 16'b0000000000000000;
		15'h1ac6: char_row_bitmap <= 16'b0000000000000000;
		15'h1ac7: char_row_bitmap <= 16'b0000000000000000;
		15'h1ac8: char_row_bitmap <= 16'b0000000000000000;
		15'h1ac9: char_row_bitmap <= 16'b0000000000000000;
		15'h1aca: char_row_bitmap <= 16'b0000000000000000;
		15'h1acb: char_row_bitmap <= 16'b0000000000000000;
		15'h1acc: char_row_bitmap <= 16'b0000000000000000;
		15'h1acd: char_row_bitmap <= 16'b0000000000000000;
		15'h1ace: char_row_bitmap <= 16'b0000000000000000;
		15'h1acf: char_row_bitmap <= 16'b0000000000000000;
		15'h1ad0: char_row_bitmap <= 16'b0000000000000000;
		15'h1ad1: char_row_bitmap <= 16'b0000000000000000;
		15'h1ad2: char_row_bitmap <= 16'b0000000000000000;
		15'h1ad3: char_row_bitmap <= 16'b0000000000000000;
		15'h1ad4: char_row_bitmap <= 16'b0000000000000000;
		15'h1ad5: char_row_bitmap <= 16'b0000000000000000;
		15'h1ad6: char_row_bitmap <= 16'b0000000000000000;
		15'h1ad7: char_row_bitmap <= 16'b0000000000000000;
		15'h1ad8: char_row_bitmap <= 16'b0000000000000000;
		15'h1ad9: char_row_bitmap <= 16'b0000000000000000;
		15'h1ada: char_row_bitmap <= 16'b0000000000000000;
		15'h1adb: char_row_bitmap <= 16'b0000000000000000;
		15'h1adc: char_row_bitmap <= 16'b0000000000000000;
		15'h1add: char_row_bitmap <= 16'b0000000000000000;
		15'h1ade: char_row_bitmap <= 16'b0000000000000000;
		15'h1adf: char_row_bitmap <= 16'b0000000000000000;
		15'h1ae0: char_row_bitmap <= 16'b0000000000000000;
		15'h1ae1: char_row_bitmap <= 16'b0000000000000000;
		15'h1ae2: char_row_bitmap <= 16'b0000000000000000;
		15'h1ae3: char_row_bitmap <= 16'b0000000000000000;
		15'h1ae4: char_row_bitmap <= 16'b0000000000000000;
		15'h1ae5: char_row_bitmap <= 16'b0000000000000000;
		15'h1ae6: char_row_bitmap <= 16'b0000000000000000;
		15'h1ae7: char_row_bitmap <= 16'b0000000000000000;
		15'h1ae8: char_row_bitmap <= 16'b0000000000000000;
		15'h1ae9: char_row_bitmap <= 16'b0000000000000000;
		15'h1aea: char_row_bitmap <= 16'b0000000000000000;
		15'h1aeb: char_row_bitmap <= 16'b0000000000000000;
		15'h1aec: char_row_bitmap <= 16'b0000000000000000;
		15'h1aed: char_row_bitmap <= 16'b0000000000000000;
		15'h1aee: char_row_bitmap <= 16'b0000000000000000;
		15'h1aef: char_row_bitmap <= 16'b0000000000000000;
		15'h1af0: char_row_bitmap <= 16'b0000000000000000;
		15'h1af1: char_row_bitmap <= 16'b0000000000000000;
		15'h1af2: char_row_bitmap <= 16'b0000000000000000;
		15'h1af3: char_row_bitmap <= 16'b0000000000000000;
		15'h1af4: char_row_bitmap <= 16'b0000000000000000;
		15'h1af5: char_row_bitmap <= 16'b0000000000000000;
		15'h1af6: char_row_bitmap <= 16'b0000000000000000;
		15'h1af7: char_row_bitmap <= 16'b0000000000000000;
		15'h1af8: char_row_bitmap <= 16'b0000000000000000;
		15'h1af9: char_row_bitmap <= 16'b0000000000000000;
		15'h1afa: char_row_bitmap <= 16'b0000000000000000;
		15'h1afb: char_row_bitmap <= 16'b0000000000000000;
		15'h1afc: char_row_bitmap <= 16'b0000000000000000;
		15'h1afd: char_row_bitmap <= 16'b0000000000000000;
		15'h1afe: char_row_bitmap <= 16'b0000000000000000;
		15'h1aff: char_row_bitmap <= 16'b0000000000000000;
		15'h1b00: char_row_bitmap <= 16'b0000000000000000;
		15'h1b01: char_row_bitmap <= 16'b0000000000000000;
		15'h1b02: char_row_bitmap <= 16'b0000000000000000;
		15'h1b03: char_row_bitmap <= 16'b0000000000000000;
		15'h1b04: char_row_bitmap <= 16'b0000000000000000;
		15'h1b05: char_row_bitmap <= 16'b0000000000000000;
		15'h1b06: char_row_bitmap <= 16'b0000000000000000;
		15'h1b07: char_row_bitmap <= 16'b0000000000000000;
		15'h1b08: char_row_bitmap <= 16'b0000000000000000;
		15'h1b09: char_row_bitmap <= 16'b0000000000000000;
		15'h1b0a: char_row_bitmap <= 16'b0000000000000000;
		15'h1b0b: char_row_bitmap <= 16'b0000000000000000;
		15'h1b0c: char_row_bitmap <= 16'b0000000000000000;
		15'h1b0d: char_row_bitmap <= 16'b0000000000000000;
		15'h1b0e: char_row_bitmap <= 16'b0000000000000000;
		15'h1b0f: char_row_bitmap <= 16'b0000000000000000;
		15'h1b10: char_row_bitmap <= 16'b0000000000000000;
		15'h1b11: char_row_bitmap <= 16'b0000000000000000;
		15'h1b12: char_row_bitmap <= 16'b0000000000000000;
		15'h1b13: char_row_bitmap <= 16'b0000000000000000;
		15'h1b14: char_row_bitmap <= 16'b0000000000000000;
		15'h1b15: char_row_bitmap <= 16'b0000000000000000;
		15'h1b16: char_row_bitmap <= 16'b0000000000000000;
		15'h1b17: char_row_bitmap <= 16'b0000000000000000;
		15'h1b18: char_row_bitmap <= 16'b0000000000000000;
		15'h1b19: char_row_bitmap <= 16'b0000000000000000;
		15'h1b1a: char_row_bitmap <= 16'b0000000000000000;
		15'h1b1b: char_row_bitmap <= 16'b0000000000000000;
		15'h1b1c: char_row_bitmap <= 16'b0000000000000000;
		15'h1b1d: char_row_bitmap <= 16'b0000000000000000;
		15'h1b1e: char_row_bitmap <= 16'b0000000000000000;
		15'h1b1f: char_row_bitmap <= 16'b0000000000000000;
		15'h1b20: char_row_bitmap <= 16'b0000000000000000;
		15'h1b21: char_row_bitmap <= 16'b0000000000000000;
		15'h1b22: char_row_bitmap <= 16'b0000000000000000;
		15'h1b23: char_row_bitmap <= 16'b0000000000000000;
		15'h1b24: char_row_bitmap <= 16'b0000000000000000;
		15'h1b25: char_row_bitmap <= 16'b0000000000000000;
		15'h1b26: char_row_bitmap <= 16'b0000000000000000;
		15'h1b27: char_row_bitmap <= 16'b0000000000000000;
		15'h1b28: char_row_bitmap <= 16'b0000000000000000;
		15'h1b29: char_row_bitmap <= 16'b0000000000000000;
		15'h1b2a: char_row_bitmap <= 16'b0000000000000000;
		15'h1b2b: char_row_bitmap <= 16'b0000000000000000;
		15'h1b2c: char_row_bitmap <= 16'b0000000000000000;
		15'h1b2d: char_row_bitmap <= 16'b0000000000000000;
		15'h1b2e: char_row_bitmap <= 16'b0000000000000000;
		15'h1b2f: char_row_bitmap <= 16'b0000000000000000;
		15'h1b30: char_row_bitmap <= 16'b0000000000000000;
		15'h1b31: char_row_bitmap <= 16'b0000000000000000;
		15'h1b32: char_row_bitmap <= 16'b0000000000000000;
		15'h1b33: char_row_bitmap <= 16'b0000000000000000;
		15'h1b34: char_row_bitmap <= 16'b0000000000000000;
		15'h1b35: char_row_bitmap <= 16'b0000000000000000;
		15'h1b36: char_row_bitmap <= 16'b0000000000000000;
		15'h1b37: char_row_bitmap <= 16'b0000000000000000;
		15'h1b38: char_row_bitmap <= 16'b0000000000000000;
		15'h1b39: char_row_bitmap <= 16'b0000000000000000;
		15'h1b3a: char_row_bitmap <= 16'b0000000000000000;
		15'h1b3b: char_row_bitmap <= 16'b0000000000000000;
		15'h1b3c: char_row_bitmap <= 16'b0000000000000000;
		15'h1b3d: char_row_bitmap <= 16'b0000000000000000;
		15'h1b3e: char_row_bitmap <= 16'b0000000000000000;
		15'h1b3f: char_row_bitmap <= 16'b0000000000000000;
		15'h1b40: char_row_bitmap <= 16'b0000000000000000;
		15'h1b41: char_row_bitmap <= 16'b0000000000000000;
		15'h1b42: char_row_bitmap <= 16'b0000000000000000;
		15'h1b43: char_row_bitmap <= 16'b0000000000000000;
		15'h1b44: char_row_bitmap <= 16'b0000000000000000;
		15'h1b45: char_row_bitmap <= 16'b0000000000000000;
		15'h1b46: char_row_bitmap <= 16'b0000000000000000;
		15'h1b47: char_row_bitmap <= 16'b0000000000000000;
		15'h1b48: char_row_bitmap <= 16'b0000000000000000;
		15'h1b49: char_row_bitmap <= 16'b0000000000000000;
		15'h1b4a: char_row_bitmap <= 16'b0000000000000000;
		15'h1b4b: char_row_bitmap <= 16'b0000000000000000;
		15'h1b4c: char_row_bitmap <= 16'b0000000000000000;
		15'h1b4d: char_row_bitmap <= 16'b0000000000000000;
		15'h1b4e: char_row_bitmap <= 16'b0000000000000000;
		15'h1b4f: char_row_bitmap <= 16'b0000000000000000;
		15'h1b50: char_row_bitmap <= 16'b0000000000000000;
		15'h1b51: char_row_bitmap <= 16'b0000000000000000;
		15'h1b52: char_row_bitmap <= 16'b0000000000000000;
		15'h1b53: char_row_bitmap <= 16'b0000000000000000;
		15'h1b54: char_row_bitmap <= 16'b0000000000000000;
		15'h1b55: char_row_bitmap <= 16'b0000000000000000;
		15'h1b56: char_row_bitmap <= 16'b0000000000000000;
		15'h1b57: char_row_bitmap <= 16'b0000000000000000;
		15'h1b58: char_row_bitmap <= 16'b0000000000000000;
		15'h1b59: char_row_bitmap <= 16'b0000000000000000;
		15'h1b5a: char_row_bitmap <= 16'b0000000000000000;
		15'h1b5b: char_row_bitmap <= 16'b0000000000000000;
		15'h1b5c: char_row_bitmap <= 16'b0000000000000000;
		15'h1b5d: char_row_bitmap <= 16'b0000000000000000;
		15'h1b5e: char_row_bitmap <= 16'b0000000000000000;
		15'h1b5f: char_row_bitmap <= 16'b0000000000000000;
		15'h1b60: char_row_bitmap <= 16'b0000000000000000;
		15'h1b61: char_row_bitmap <= 16'b0000000000000000;
		15'h1b62: char_row_bitmap <= 16'b0000000000000000;
		15'h1b63: char_row_bitmap <= 16'b0000000000000000;
		15'h1b64: char_row_bitmap <= 16'b0000000000000000;
		15'h1b65: char_row_bitmap <= 16'b0000000000000000;
		15'h1b66: char_row_bitmap <= 16'b0000000000000000;
		15'h1b67: char_row_bitmap <= 16'b0000000000000000;
		15'h1b68: char_row_bitmap <= 16'b0000000000000000;
		15'h1b69: char_row_bitmap <= 16'b0000000000000000;
		15'h1b6a: char_row_bitmap <= 16'b0000000000000000;
		15'h1b6b: char_row_bitmap <= 16'b0000000000000000;
		15'h1b6c: char_row_bitmap <= 16'b0000000000000000;
		15'h1b6d: char_row_bitmap <= 16'b0000000000000000;
		15'h1b6e: char_row_bitmap <= 16'b0000000000000000;
		15'h1b6f: char_row_bitmap <= 16'b0000000000000000;
		15'h1b70: char_row_bitmap <= 16'b0000000000000000;
		15'h1b71: char_row_bitmap <= 16'b0000000000000000;
		15'h1b72: char_row_bitmap <= 16'b0000000000000000;
		15'h1b73: char_row_bitmap <= 16'b0000000000000000;
		15'h1b74: char_row_bitmap <= 16'b0000000000000000;
		15'h1b75: char_row_bitmap <= 16'b0000000000000000;
		15'h1b76: char_row_bitmap <= 16'b0000000000000000;
		15'h1b77: char_row_bitmap <= 16'b0000000000000000;
		15'h1b78: char_row_bitmap <= 16'b0000000000000000;
		15'h1b79: char_row_bitmap <= 16'b0000000000000000;
		15'h1b7a: char_row_bitmap <= 16'b0000000000000000;
		15'h1b7b: char_row_bitmap <= 16'b0000000000000000;
		15'h1b7c: char_row_bitmap <= 16'b0000000000000000;
		15'h1b7d: char_row_bitmap <= 16'b0000000000000000;
		15'h1b7e: char_row_bitmap <= 16'b0000000000000000;
		15'h1b7f: char_row_bitmap <= 16'b0000000000000000;
		15'h1b80: char_row_bitmap <= 16'b0000000000000000;
		15'h1b81: char_row_bitmap <= 16'b0000000000000000;
		15'h1b82: char_row_bitmap <= 16'b0000000000000000;
		15'h1b83: char_row_bitmap <= 16'b0000000000000000;
		15'h1b84: char_row_bitmap <= 16'b0000000000000000;
		15'h1b85: char_row_bitmap <= 16'b0000000000000000;
		15'h1b86: char_row_bitmap <= 16'b0000000000000000;
		15'h1b87: char_row_bitmap <= 16'b0000000000000000;
		15'h1b88: char_row_bitmap <= 16'b0000000000000000;
		15'h1b89: char_row_bitmap <= 16'b0000000000000000;
		15'h1b8a: char_row_bitmap <= 16'b0000000000000000;
		15'h1b8b: char_row_bitmap <= 16'b0000000000000000;
		15'h1b8c: char_row_bitmap <= 16'b0000000000000000;
		15'h1b8d: char_row_bitmap <= 16'b0000000000000000;
		15'h1b8e: char_row_bitmap <= 16'b0000000000000000;
		15'h1b8f: char_row_bitmap <= 16'b0000000000000000;
		15'h1b90: char_row_bitmap <= 16'b0000000000000000;
		15'h1b91: char_row_bitmap <= 16'b0000000000000000;
		15'h1b92: char_row_bitmap <= 16'b0000000000000000;
		15'h1b93: char_row_bitmap <= 16'b0000000000000000;
		15'h1b94: char_row_bitmap <= 16'b0000000000000000;
		15'h1b95: char_row_bitmap <= 16'b0000000000000000;
		15'h1b96: char_row_bitmap <= 16'b0000000000000000;
		15'h1b97: char_row_bitmap <= 16'b0000000000000000;
		15'h1b98: char_row_bitmap <= 16'b0000000000000000;
		15'h1b99: char_row_bitmap <= 16'b0000000000000000;
		15'h1b9a: char_row_bitmap <= 16'b0000000000000000;
		15'h1b9b: char_row_bitmap <= 16'b0000000000000000;
		15'h1b9c: char_row_bitmap <= 16'b0000000000000000;
		15'h1b9d: char_row_bitmap <= 16'b0000000000000000;
		15'h1b9e: char_row_bitmap <= 16'b0000000000000000;
		15'h1b9f: char_row_bitmap <= 16'b0000000000000000;
		15'h1ba0: char_row_bitmap <= 16'b0000000000000000;
		15'h1ba1: char_row_bitmap <= 16'b0000000000000000;
		15'h1ba2: char_row_bitmap <= 16'b0000000000000000;
		15'h1ba3: char_row_bitmap <= 16'b0000000000000000;
		15'h1ba4: char_row_bitmap <= 16'b0000000000000000;
		15'h1ba5: char_row_bitmap <= 16'b0000000000000000;
		15'h1ba6: char_row_bitmap <= 16'b0000000000000000;
		15'h1ba7: char_row_bitmap <= 16'b0000000000000000;
		15'h1ba8: char_row_bitmap <= 16'b0000000000000000;
		15'h1ba9: char_row_bitmap <= 16'b0000000000000000;
		15'h1baa: char_row_bitmap <= 16'b0000000000000000;
		15'h1bab: char_row_bitmap <= 16'b0000000000000000;
		15'h1bac: char_row_bitmap <= 16'b0000000000000000;
		15'h1bad: char_row_bitmap <= 16'b0000000000000000;
		15'h1bae: char_row_bitmap <= 16'b0000000000000000;
		15'h1baf: char_row_bitmap <= 16'b0000000000000000;
		15'h1bb0: char_row_bitmap <= 16'b0000000000000000;
		15'h1bb1: char_row_bitmap <= 16'b0000000000000000;
		15'h1bb2: char_row_bitmap <= 16'b0000000000000000;
		15'h1bb3: char_row_bitmap <= 16'b0000000000000000;
		15'h1bb4: char_row_bitmap <= 16'b0000000000000000;
		15'h1bb5: char_row_bitmap <= 16'b0000000000000000;
		15'h1bb6: char_row_bitmap <= 16'b0000000000000000;
		15'h1bb7: char_row_bitmap <= 16'b0000000000000000;
		15'h1bb8: char_row_bitmap <= 16'b0000000000000000;
		15'h1bb9: char_row_bitmap <= 16'b0000000000000000;
		15'h1bba: char_row_bitmap <= 16'b0000000000000000;
		15'h1bbb: char_row_bitmap <= 16'b0000000000000000;
		15'h1bbc: char_row_bitmap <= 16'b0000000000000000;
		15'h1bbd: char_row_bitmap <= 16'b0000000000000000;
		15'h1bbe: char_row_bitmap <= 16'b0000000000000000;
		15'h1bbf: char_row_bitmap <= 16'b0000000000000000;
		15'h1bc0: char_row_bitmap <= 16'b0000000000000000;
		15'h1bc1: char_row_bitmap <= 16'b0000000000000000;
		15'h1bc2: char_row_bitmap <= 16'b0000000000000000;
		15'h1bc3: char_row_bitmap <= 16'b0000000000000000;
		15'h1bc4: char_row_bitmap <= 16'b0000000000000000;
		15'h1bc5: char_row_bitmap <= 16'b0000000000000000;
		15'h1bc6: char_row_bitmap <= 16'b0000000000000000;
		15'h1bc7: char_row_bitmap <= 16'b0000000000000000;
		15'h1bc8: char_row_bitmap <= 16'b0000000000000000;
		15'h1bc9: char_row_bitmap <= 16'b0000000000000000;
		15'h1bca: char_row_bitmap <= 16'b0000000000000000;
		15'h1bcb: char_row_bitmap <= 16'b0000000000000000;
		15'h1bcc: char_row_bitmap <= 16'b0000000000000000;
		15'h1bcd: char_row_bitmap <= 16'b0000000000000000;
		15'h1bce: char_row_bitmap <= 16'b0000000000000000;
		15'h1bcf: char_row_bitmap <= 16'b0000000000000000;
		15'h1bd0: char_row_bitmap <= 16'b0000000000000000;
		15'h1bd1: char_row_bitmap <= 16'b0000000000000000;
		15'h1bd2: char_row_bitmap <= 16'b0000000000000000;
		15'h1bd3: char_row_bitmap <= 16'b0000000000000000;
		15'h1bd4: char_row_bitmap <= 16'b0000000000000000;
		15'h1bd5: char_row_bitmap <= 16'b0000000000000000;
		15'h1bd6: char_row_bitmap <= 16'b0000000000000000;
		15'h1bd7: char_row_bitmap <= 16'b0000000000000000;
		15'h1bd8: char_row_bitmap <= 16'b0000000000000000;
		15'h1bd9: char_row_bitmap <= 16'b0000000000000000;
		15'h1bda: char_row_bitmap <= 16'b0000000000000000;
		15'h1bdb: char_row_bitmap <= 16'b0000000000000000;
		15'h1bdc: char_row_bitmap <= 16'b0000000000000000;
		15'h1bdd: char_row_bitmap <= 16'b0000000000000000;
		15'h1bde: char_row_bitmap <= 16'b0000000000000000;
		15'h1bdf: char_row_bitmap <= 16'b0000000000000000;
		15'h1be0: char_row_bitmap <= 16'b0000000000000000;
		15'h1be1: char_row_bitmap <= 16'b0000000000000000;
		15'h1be2: char_row_bitmap <= 16'b0000000000000000;
		15'h1be3: char_row_bitmap <= 16'b0000000000000000;
		15'h1be4: char_row_bitmap <= 16'b0000000000000000;
		15'h1be5: char_row_bitmap <= 16'b0000000000000000;
		15'h1be6: char_row_bitmap <= 16'b0000000000000000;
		15'h1be7: char_row_bitmap <= 16'b0000000000000000;
		15'h1be8: char_row_bitmap <= 16'b0000000000000000;
		15'h1be9: char_row_bitmap <= 16'b0000000000000000;
		15'h1bea: char_row_bitmap <= 16'b0000000000000000;
		15'h1beb: char_row_bitmap <= 16'b0000000000000000;
		15'h1bec: char_row_bitmap <= 16'b0000000000000000;
		15'h1bed: char_row_bitmap <= 16'b0000000000000000;
		15'h1bee: char_row_bitmap <= 16'b0000000000000000;
		15'h1bef: char_row_bitmap <= 16'b0000000000000000;
		15'h1bf0: char_row_bitmap <= 16'b0000000000000000;
		15'h1bf1: char_row_bitmap <= 16'b0000000000000000;
		15'h1bf2: char_row_bitmap <= 16'b0000000000000000;
		15'h1bf3: char_row_bitmap <= 16'b0000000000000000;
		15'h1bf4: char_row_bitmap <= 16'b0000000000000000;
		15'h1bf5: char_row_bitmap <= 16'b0000000000000000;
		15'h1bf6: char_row_bitmap <= 16'b0000000000000000;
		15'h1bf7: char_row_bitmap <= 16'b0000000000000000;
		15'h1bf8: char_row_bitmap <= 16'b0000000000000000;
		15'h1bf9: char_row_bitmap <= 16'b0000000000000000;
		15'h1bfa: char_row_bitmap <= 16'b0000000000000000;
		15'h1bfb: char_row_bitmap <= 16'b0000000000000000;
		15'h1bfc: char_row_bitmap <= 16'b0000000000000000;
		15'h1bfd: char_row_bitmap <= 16'b0000000000000000;
		15'h1bfe: char_row_bitmap <= 16'b0000000000000000;
		15'h1bff: char_row_bitmap <= 16'b0000000000000000;
		15'h1c00: char_row_bitmap <= 16'b0000000000000000;
		15'h1c01: char_row_bitmap <= 16'b0000000000000000;
		15'h1c02: char_row_bitmap <= 16'b0000000000000000;
		15'h1c03: char_row_bitmap <= 16'b0000000000000000;
		15'h1c04: char_row_bitmap <= 16'b0000000000000000;
		15'h1c05: char_row_bitmap <= 16'b0000000000000000;
		15'h1c06: char_row_bitmap <= 16'b0000000000000000;
		15'h1c07: char_row_bitmap <= 16'b0000000000000000;
		15'h1c08: char_row_bitmap <= 16'b0000000000000000;
		15'h1c09: char_row_bitmap <= 16'b0000000000000000;
		15'h1c0a: char_row_bitmap <= 16'b0000000000000000;
		15'h1c0b: char_row_bitmap <= 16'b0000000000000000;
		15'h1c0c: char_row_bitmap <= 16'b0000000000000000;
		15'h1c0d: char_row_bitmap <= 16'b0000000000000000;
		15'h1c0e: char_row_bitmap <= 16'b0000000000000000;
		15'h1c0f: char_row_bitmap <= 16'b0000000000000000;
		15'h1c10: char_row_bitmap <= 16'b0000000000000000;
		15'h1c11: char_row_bitmap <= 16'b0000000000000000;
		15'h1c12: char_row_bitmap <= 16'b0000000000000000;
		15'h1c13: char_row_bitmap <= 16'b0000000000000000;
		15'h1c14: char_row_bitmap <= 16'b0000000000000000;
		15'h1c15: char_row_bitmap <= 16'b0000000000000000;
		15'h1c16: char_row_bitmap <= 16'b0000000000000000;
		15'h1c17: char_row_bitmap <= 16'b0000000000000000;
		15'h1c18: char_row_bitmap <= 16'b0000000000000000;
		15'h1c19: char_row_bitmap <= 16'b0000000000000000;
		15'h1c1a: char_row_bitmap <= 16'b0000000000000000;
		15'h1c1b: char_row_bitmap <= 16'b0000000000000000;
		15'h1c1c: char_row_bitmap <= 16'b0000000000000000;
		15'h1c1d: char_row_bitmap <= 16'b0000000000000000;
		15'h1c1e: char_row_bitmap <= 16'b0000000000000000;
		15'h1c1f: char_row_bitmap <= 16'b0000000000000000;
		15'h1c20: char_row_bitmap <= 16'b0000000000000000;
		15'h1c21: char_row_bitmap <= 16'b0000000000000000;
		15'h1c22: char_row_bitmap <= 16'b0000000000000000;
		15'h1c23: char_row_bitmap <= 16'b0000000000000000;
		15'h1c24: char_row_bitmap <= 16'b0000000000000000;
		15'h1c25: char_row_bitmap <= 16'b0000000000000000;
		15'h1c26: char_row_bitmap <= 16'b0000000000000000;
		15'h1c27: char_row_bitmap <= 16'b0000000000000000;
		15'h1c28: char_row_bitmap <= 16'b0000000000000000;
		15'h1c29: char_row_bitmap <= 16'b0000000000000000;
		15'h1c2a: char_row_bitmap <= 16'b0000000000000000;
		15'h1c2b: char_row_bitmap <= 16'b0000000000000000;
		15'h1c2c: char_row_bitmap <= 16'b0000000000000000;
		15'h1c2d: char_row_bitmap <= 16'b0000000000000000;
		15'h1c2e: char_row_bitmap <= 16'b0000000000000000;
		15'h1c2f: char_row_bitmap <= 16'b0000000000000000;
		15'h1c30: char_row_bitmap <= 16'b0000000000000000;
		15'h1c31: char_row_bitmap <= 16'b0000000000000000;
		15'h1c32: char_row_bitmap <= 16'b0000000000000000;
		15'h1c33: char_row_bitmap <= 16'b0000000000000000;
		15'h1c34: char_row_bitmap <= 16'b0000000000000000;
		15'h1c35: char_row_bitmap <= 16'b0000000000000000;
		15'h1c36: char_row_bitmap <= 16'b0000000000000000;
		15'h1c37: char_row_bitmap <= 16'b0000000000000000;
		15'h1c38: char_row_bitmap <= 16'b0000000000000000;
		15'h1c39: char_row_bitmap <= 16'b0000000000000000;
		15'h1c3a: char_row_bitmap <= 16'b0000000000000000;
		15'h1c3b: char_row_bitmap <= 16'b0000000000000000;
		15'h1c3c: char_row_bitmap <= 16'b0000000000000000;
		15'h1c3d: char_row_bitmap <= 16'b0000000000000000;
		15'h1c3e: char_row_bitmap <= 16'b0000000000000000;
		15'h1c3f: char_row_bitmap <= 16'b0000000000000000;
		15'h1c40: char_row_bitmap <= 16'b0000000000000000;
		15'h1c41: char_row_bitmap <= 16'b0000000000000000;
		15'h1c42: char_row_bitmap <= 16'b0000000000000000;
		15'h1c43: char_row_bitmap <= 16'b0000000000000000;
		15'h1c44: char_row_bitmap <= 16'b0000000000000000;
		15'h1c45: char_row_bitmap <= 16'b0000000000000000;
		15'h1c46: char_row_bitmap <= 16'b0000000000000000;
		15'h1c47: char_row_bitmap <= 16'b0000000000000000;
		15'h1c48: char_row_bitmap <= 16'b0000000000000000;
		15'h1c49: char_row_bitmap <= 16'b0000000000000000;
		15'h1c4a: char_row_bitmap <= 16'b0000000000000000;
		15'h1c4b: char_row_bitmap <= 16'b0000000000000000;
		15'h1c4c: char_row_bitmap <= 16'b0000000000000000;
		15'h1c4d: char_row_bitmap <= 16'b0000000000000000;
		15'h1c4e: char_row_bitmap <= 16'b0000000000000000;
		15'h1c4f: char_row_bitmap <= 16'b0000000000000000;
		15'h1c50: char_row_bitmap <= 16'b0000000000000000;
		15'h1c51: char_row_bitmap <= 16'b0000000000000000;
		15'h1c52: char_row_bitmap <= 16'b0000000000000000;
		15'h1c53: char_row_bitmap <= 16'b0000000000000000;
		15'h1c54: char_row_bitmap <= 16'b0000000000000000;
		15'h1c55: char_row_bitmap <= 16'b0000000000000000;
		15'h1c56: char_row_bitmap <= 16'b0000000000000000;
		15'h1c57: char_row_bitmap <= 16'b0000000000000000;
		15'h1c58: char_row_bitmap <= 16'b0000000000000000;
		15'h1c59: char_row_bitmap <= 16'b0000000000000000;
		15'h1c5a: char_row_bitmap <= 16'b0000000000000000;
		15'h1c5b: char_row_bitmap <= 16'b0000000000000000;
		15'h1c5c: char_row_bitmap <= 16'b0000000000000000;
		15'h1c5d: char_row_bitmap <= 16'b0000000000000000;
		15'h1c5e: char_row_bitmap <= 16'b0000000000000000;
		15'h1c5f: char_row_bitmap <= 16'b0000000000000000;
		15'h1c60: char_row_bitmap <= 16'b0000000000000000;
		15'h1c61: char_row_bitmap <= 16'b0000000000000000;
		15'h1c62: char_row_bitmap <= 16'b0000000000000000;
		15'h1c63: char_row_bitmap <= 16'b0000000000000000;
		15'h1c64: char_row_bitmap <= 16'b0000000000000000;
		15'h1c65: char_row_bitmap <= 16'b0000000000000000;
		15'h1c66: char_row_bitmap <= 16'b0000000000000000;
		15'h1c67: char_row_bitmap <= 16'b0000000000000000;
		15'h1c68: char_row_bitmap <= 16'b0000000000000000;
		15'h1c69: char_row_bitmap <= 16'b0000000000000000;
		15'h1c6a: char_row_bitmap <= 16'b0000000000000000;
		15'h1c6b: char_row_bitmap <= 16'b0000000000000000;
		15'h1c6c: char_row_bitmap <= 16'b0000000000000000;
		15'h1c6d: char_row_bitmap <= 16'b0000000000000000;
		15'h1c6e: char_row_bitmap <= 16'b0000000000000000;
		15'h1c6f: char_row_bitmap <= 16'b0000000000000000;
		15'h1c70: char_row_bitmap <= 16'b0000000000000000;
		15'h1c71: char_row_bitmap <= 16'b0000000000000000;
		15'h1c72: char_row_bitmap <= 16'b0000000000000000;
		15'h1c73: char_row_bitmap <= 16'b0000000000000000;
		15'h1c74: char_row_bitmap <= 16'b0000000000000000;
		15'h1c75: char_row_bitmap <= 16'b0000000000000000;
		15'h1c76: char_row_bitmap <= 16'b0000000000000000;
		15'h1c77: char_row_bitmap <= 16'b0000000000000000;
		15'h1c78: char_row_bitmap <= 16'b0000000000000000;
		15'h1c79: char_row_bitmap <= 16'b0000000000000000;
		15'h1c7a: char_row_bitmap <= 16'b0000000000000000;
		15'h1c7b: char_row_bitmap <= 16'b0000000000000000;
		15'h1c7c: char_row_bitmap <= 16'b0000000000000000;
		15'h1c7d: char_row_bitmap <= 16'b0000000000000000;
		15'h1c7e: char_row_bitmap <= 16'b0000000000000000;
		15'h1c7f: char_row_bitmap <= 16'b0000000000000000;
		15'h1c80: char_row_bitmap <= 16'b0000000000000000;
		15'h1c81: char_row_bitmap <= 16'b0000000000000000;
		15'h1c82: char_row_bitmap <= 16'b0000000000000000;
		15'h1c83: char_row_bitmap <= 16'b0000000000000000;
		15'h1c84: char_row_bitmap <= 16'b0000000000000000;
		15'h1c85: char_row_bitmap <= 16'b0000000000000000;
		15'h1c86: char_row_bitmap <= 16'b0000000000000000;
		15'h1c87: char_row_bitmap <= 16'b0000000000000000;
		15'h1c88: char_row_bitmap <= 16'b0000000000000000;
		15'h1c89: char_row_bitmap <= 16'b0000000000000000;
		15'h1c8a: char_row_bitmap <= 16'b0000000000000000;
		15'h1c8b: char_row_bitmap <= 16'b0000000000000000;
		15'h1c8c: char_row_bitmap <= 16'b0000000000000000;
		15'h1c8d: char_row_bitmap <= 16'b0000000000000000;
		15'h1c8e: char_row_bitmap <= 16'b0000000000000000;
		15'h1c8f: char_row_bitmap <= 16'b0000000000000000;
		15'h1c90: char_row_bitmap <= 16'b0000000000000000;
		15'h1c91: char_row_bitmap <= 16'b0000000000000000;
		15'h1c92: char_row_bitmap <= 16'b0000000000000000;
		15'h1c93: char_row_bitmap <= 16'b0000000000000000;
		15'h1c94: char_row_bitmap <= 16'b0000000000000000;
		15'h1c95: char_row_bitmap <= 16'b0000000000000000;
		15'h1c96: char_row_bitmap <= 16'b0000000000000000;
		15'h1c97: char_row_bitmap <= 16'b0000000000000000;
		15'h1c98: char_row_bitmap <= 16'b0000000000000000;
		15'h1c99: char_row_bitmap <= 16'b0000000000000000;
		15'h1c9a: char_row_bitmap <= 16'b0000000000000000;
		15'h1c9b: char_row_bitmap <= 16'b0000000000000000;
		15'h1c9c: char_row_bitmap <= 16'b0000000000000000;
		15'h1c9d: char_row_bitmap <= 16'b0000000000000000;
		15'h1c9e: char_row_bitmap <= 16'b0000000000000000;
		15'h1c9f: char_row_bitmap <= 16'b0000000000000000;
		15'h1ca0: char_row_bitmap <= 16'b0000000000000000;
		15'h1ca1: char_row_bitmap <= 16'b0000000000000000;
		15'h1ca2: char_row_bitmap <= 16'b0000000000000000;
		15'h1ca3: char_row_bitmap <= 16'b0000000000000000;
		15'h1ca4: char_row_bitmap <= 16'b0000000000000000;
		15'h1ca5: char_row_bitmap <= 16'b0000000000000000;
		15'h1ca6: char_row_bitmap <= 16'b0000000000000000;
		15'h1ca7: char_row_bitmap <= 16'b0000000000000000;
		15'h1ca8: char_row_bitmap <= 16'b0000000000000000;
		15'h1ca9: char_row_bitmap <= 16'b0000000000000000;
		15'h1caa: char_row_bitmap <= 16'b0000000000000000;
		15'h1cab: char_row_bitmap <= 16'b0000000000000000;
		15'h1cac: char_row_bitmap <= 16'b0000000000000000;
		15'h1cad: char_row_bitmap <= 16'b0000000000000000;
		15'h1cae: char_row_bitmap <= 16'b0000000000000000;
		15'h1caf: char_row_bitmap <= 16'b0000000000000000;
		15'h1cb0: char_row_bitmap <= 16'b0000000000000000;
		15'h1cb1: char_row_bitmap <= 16'b0000000000000000;
		15'h1cb2: char_row_bitmap <= 16'b0000000000000000;
		15'h1cb3: char_row_bitmap <= 16'b0000000000000000;
		15'h1cb4: char_row_bitmap <= 16'b0000000000000000;
		15'h1cb5: char_row_bitmap <= 16'b0000000000000000;
		15'h1cb6: char_row_bitmap <= 16'b0000000000000000;
		15'h1cb7: char_row_bitmap <= 16'b0000000000000000;
		15'h1cb8: char_row_bitmap <= 16'b0000000000000000;
		15'h1cb9: char_row_bitmap <= 16'b0000000000000000;
		15'h1cba: char_row_bitmap <= 16'b0000000000000000;
		15'h1cbb: char_row_bitmap <= 16'b0000000000000000;
		15'h1cbc: char_row_bitmap <= 16'b0000000000000000;
		15'h1cbd: char_row_bitmap <= 16'b0000000000000000;
		15'h1cbe: char_row_bitmap <= 16'b0000000000000000;
		15'h1cbf: char_row_bitmap <= 16'b0000000000000000;
		15'h1cc0: char_row_bitmap <= 16'b0000000000000000;
		15'h1cc1: char_row_bitmap <= 16'b0000000000000000;
		15'h1cc2: char_row_bitmap <= 16'b0000000000000000;
		15'h1cc3: char_row_bitmap <= 16'b0000000000000000;
		15'h1cc4: char_row_bitmap <= 16'b0000000000000000;
		15'h1cc5: char_row_bitmap <= 16'b0000000000000000;
		15'h1cc6: char_row_bitmap <= 16'b0000000000000000;
		15'h1cc7: char_row_bitmap <= 16'b0000000000000000;
		15'h1cc8: char_row_bitmap <= 16'b0000000000000000;
		15'h1cc9: char_row_bitmap <= 16'b0000000000000000;
		15'h1cca: char_row_bitmap <= 16'b0000000000000000;
		15'h1ccb: char_row_bitmap <= 16'b0000000000000000;
		15'h1ccc: char_row_bitmap <= 16'b0000000000000000;
		15'h1ccd: char_row_bitmap <= 16'b0000000000000000;
		15'h1cce: char_row_bitmap <= 16'b0000000000000000;
		15'h1ccf: char_row_bitmap <= 16'b0000000000000000;
		15'h1cd0: char_row_bitmap <= 16'b0000000000000000;
		15'h1cd1: char_row_bitmap <= 16'b0000000000000000;
		15'h1cd2: char_row_bitmap <= 16'b0000000000000000;
		15'h1cd3: char_row_bitmap <= 16'b0000000000000000;
		15'h1cd4: char_row_bitmap <= 16'b0000000000000000;
		15'h1cd5: char_row_bitmap <= 16'b0000000000000000;
		15'h1cd6: char_row_bitmap <= 16'b0000000000000000;
		15'h1cd7: char_row_bitmap <= 16'b0000000000000000;
		15'h1cd8: char_row_bitmap <= 16'b0000000000000000;
		15'h1cd9: char_row_bitmap <= 16'b0000000000000000;
		15'h1cda: char_row_bitmap <= 16'b0000000000000000;
		15'h1cdb: char_row_bitmap <= 16'b0000000000000000;
		15'h1cdc: char_row_bitmap <= 16'b0000000000000000;
		15'h1cdd: char_row_bitmap <= 16'b0000000000000000;
		15'h1cde: char_row_bitmap <= 16'b0000000000000000;
		15'h1cdf: char_row_bitmap <= 16'b0000000000000000;
		15'h1ce0: char_row_bitmap <= 16'b0000000000000000;
		15'h1ce1: char_row_bitmap <= 16'b0000000000000000;
		15'h1ce2: char_row_bitmap <= 16'b0000000000000000;
		15'h1ce3: char_row_bitmap <= 16'b0000000000000000;
		15'h1ce4: char_row_bitmap <= 16'b0000000000000000;
		15'h1ce5: char_row_bitmap <= 16'b0000000000000000;
		15'h1ce6: char_row_bitmap <= 16'b0000000000000000;
		15'h1ce7: char_row_bitmap <= 16'b0000000000000000;
		15'h1ce8: char_row_bitmap <= 16'b0000000000000000;
		15'h1ce9: char_row_bitmap <= 16'b0000000000000000;
		15'h1cea: char_row_bitmap <= 16'b0000000000000000;
		15'h1ceb: char_row_bitmap <= 16'b0000000000000000;
		15'h1cec: char_row_bitmap <= 16'b0000000000000000;
		15'h1ced: char_row_bitmap <= 16'b0000000000000000;
		15'h1cee: char_row_bitmap <= 16'b0000000000000000;
		15'h1cef: char_row_bitmap <= 16'b0000000000000000;
		15'h1cf0: char_row_bitmap <= 16'b0000000000000000;
		15'h1cf1: char_row_bitmap <= 16'b0000000000000000;
		15'h1cf2: char_row_bitmap <= 16'b0000000000000000;
		15'h1cf3: char_row_bitmap <= 16'b0000000000000000;
		15'h1cf4: char_row_bitmap <= 16'b0000000000000000;
		15'h1cf5: char_row_bitmap <= 16'b0000000000000000;
		15'h1cf6: char_row_bitmap <= 16'b0000000000000000;
		15'h1cf7: char_row_bitmap <= 16'b0000000000000000;
		15'h1cf8: char_row_bitmap <= 16'b0000000000000000;
		15'h1cf9: char_row_bitmap <= 16'b0000000000000000;
		15'h1cfa: char_row_bitmap <= 16'b0000000000000000;
		15'h1cfb: char_row_bitmap <= 16'b0000000000000000;
		15'h1cfc: char_row_bitmap <= 16'b0000000000000000;
		15'h1cfd: char_row_bitmap <= 16'b0000000000000000;
		15'h1cfe: char_row_bitmap <= 16'b0000000000000000;
		15'h1cff: char_row_bitmap <= 16'b0000000000000000;
		15'h1d00: char_row_bitmap <= 16'b0000000000000000;
		15'h1d01: char_row_bitmap <= 16'b0000000000000000;
		15'h1d02: char_row_bitmap <= 16'b0000000000000000;
		15'h1d03: char_row_bitmap <= 16'b0000000000000000;
		15'h1d04: char_row_bitmap <= 16'b0000000000000000;
		15'h1d05: char_row_bitmap <= 16'b0000000000000000;
		15'h1d06: char_row_bitmap <= 16'b0000000000000000;
		15'h1d07: char_row_bitmap <= 16'b0000000000000000;
		15'h1d08: char_row_bitmap <= 16'b0000000000000000;
		15'h1d09: char_row_bitmap <= 16'b0000000000000000;
		15'h1d0a: char_row_bitmap <= 16'b0000000000000000;
		15'h1d0b: char_row_bitmap <= 16'b0000000000000000;
		15'h1d0c: char_row_bitmap <= 16'b0000000000000000;
		15'h1d0d: char_row_bitmap <= 16'b0000000000000000;
		15'h1d0e: char_row_bitmap <= 16'b0000000000000000;
		15'h1d0f: char_row_bitmap <= 16'b0000000000000000;
		15'h1d10: char_row_bitmap <= 16'b0000000000000000;
		15'h1d11: char_row_bitmap <= 16'b0000000000000000;
		15'h1d12: char_row_bitmap <= 16'b0000000000000000;
		15'h1d13: char_row_bitmap <= 16'b0000000000000000;
		15'h1d14: char_row_bitmap <= 16'b0000000000000000;
		15'h1d15: char_row_bitmap <= 16'b0000000000000000;
		15'h1d16: char_row_bitmap <= 16'b0000000000000000;
		15'h1d17: char_row_bitmap <= 16'b0000000000000000;
		15'h1d18: char_row_bitmap <= 16'b0000000000000000;
		15'h1d19: char_row_bitmap <= 16'b0000000000000000;
		15'h1d1a: char_row_bitmap <= 16'b0000000000000000;
		15'h1d1b: char_row_bitmap <= 16'b0000000000000000;
		15'h1d1c: char_row_bitmap <= 16'b0000000000000000;
		15'h1d1d: char_row_bitmap <= 16'b0000000000000000;
		15'h1d1e: char_row_bitmap <= 16'b0000000000000000;
		15'h1d1f: char_row_bitmap <= 16'b0000000000000000;
		15'h1d20: char_row_bitmap <= 16'b0000000000000000;
		15'h1d21: char_row_bitmap <= 16'b0000000000000000;
		15'h1d22: char_row_bitmap <= 16'b0000000000000000;
		15'h1d23: char_row_bitmap <= 16'b0000000000000000;
		15'h1d24: char_row_bitmap <= 16'b0000000000000000;
		15'h1d25: char_row_bitmap <= 16'b0000000000000000;
		15'h1d26: char_row_bitmap <= 16'b0000000000000000;
		15'h1d27: char_row_bitmap <= 16'b0000000000000000;
		15'h1d28: char_row_bitmap <= 16'b0000000000000000;
		15'h1d29: char_row_bitmap <= 16'b0000000000000000;
		15'h1d2a: char_row_bitmap <= 16'b0000000000000000;
		15'h1d2b: char_row_bitmap <= 16'b0000000000000000;
		15'h1d2c: char_row_bitmap <= 16'b0000000000000000;
		15'h1d2d: char_row_bitmap <= 16'b0000000000000000;
		15'h1d2e: char_row_bitmap <= 16'b0000000000000000;
		15'h1d2f: char_row_bitmap <= 16'b0000000000000000;
		15'h1d30: char_row_bitmap <= 16'b0000000000000000;
		15'h1d31: char_row_bitmap <= 16'b0000000000000000;
		15'h1d32: char_row_bitmap <= 16'b0000000000000000;
		15'h1d33: char_row_bitmap <= 16'b0000000000000000;
		15'h1d34: char_row_bitmap <= 16'b0000000000000000;
		15'h1d35: char_row_bitmap <= 16'b0000000000000000;
		15'h1d36: char_row_bitmap <= 16'b0000000000000000;
		15'h1d37: char_row_bitmap <= 16'b0000000000000000;
		15'h1d38: char_row_bitmap <= 16'b0000000000000000;
		15'h1d39: char_row_bitmap <= 16'b0000000000000000;
		15'h1d3a: char_row_bitmap <= 16'b0000000000000000;
		15'h1d3b: char_row_bitmap <= 16'b0000000000000000;
		15'h1d3c: char_row_bitmap <= 16'b0000000000000000;
		15'h1d3d: char_row_bitmap <= 16'b0000000000000000;
		15'h1d3e: char_row_bitmap <= 16'b0000000000000000;
		15'h1d3f: char_row_bitmap <= 16'b0000000000000000;
		15'h1d40: char_row_bitmap <= 16'b0000000000000000;
		15'h1d41: char_row_bitmap <= 16'b0000000000000000;
		15'h1d42: char_row_bitmap <= 16'b0000000000000000;
		15'h1d43: char_row_bitmap <= 16'b0000000000000000;
		15'h1d44: char_row_bitmap <= 16'b0000000000000000;
		15'h1d45: char_row_bitmap <= 16'b0000000000000000;
		15'h1d46: char_row_bitmap <= 16'b0000000000000000;
		15'h1d47: char_row_bitmap <= 16'b0000000000000000;
		15'h1d48: char_row_bitmap <= 16'b0000000000000000;
		15'h1d49: char_row_bitmap <= 16'b0000000000000000;
		15'h1d4a: char_row_bitmap <= 16'b0000000000000000;
		15'h1d4b: char_row_bitmap <= 16'b0000000000000000;
		15'h1d4c: char_row_bitmap <= 16'b0000000000000000;
		15'h1d4d: char_row_bitmap <= 16'b0000000000000000;
		15'h1d4e: char_row_bitmap <= 16'b0000000000000000;
		15'h1d4f: char_row_bitmap <= 16'b0000000000000000;
		15'h1d50: char_row_bitmap <= 16'b0000000000000000;
		15'h1d51: char_row_bitmap <= 16'b0000000000000000;
		15'h1d52: char_row_bitmap <= 16'b0000000000000000;
		15'h1d53: char_row_bitmap <= 16'b0000000000000000;
		15'h1d54: char_row_bitmap <= 16'b0000000000000000;
		15'h1d55: char_row_bitmap <= 16'b0000000000000000;
		15'h1d56: char_row_bitmap <= 16'b0000000000000000;
		15'h1d57: char_row_bitmap <= 16'b0000000000000000;
		15'h1d58: char_row_bitmap <= 16'b0000000000000000;
		15'h1d59: char_row_bitmap <= 16'b0000000000000000;
		15'h1d5a: char_row_bitmap <= 16'b0000000000000000;
		15'h1d5b: char_row_bitmap <= 16'b0000000000000000;
		15'h1d5c: char_row_bitmap <= 16'b0000000000000000;
		15'h1d5d: char_row_bitmap <= 16'b0000000000000000;
		15'h1d5e: char_row_bitmap <= 16'b0000000000000000;
		15'h1d5f: char_row_bitmap <= 16'b0000000000000000;
		15'h1d60: char_row_bitmap <= 16'b0000000000000000;
		15'h1d61: char_row_bitmap <= 16'b0000000000000000;
		15'h1d62: char_row_bitmap <= 16'b0000000000000000;
		15'h1d63: char_row_bitmap <= 16'b0000000000000000;
		15'h1d64: char_row_bitmap <= 16'b0000000000000000;
		15'h1d65: char_row_bitmap <= 16'b0000000000000000;
		15'h1d66: char_row_bitmap <= 16'b0000000000000000;
		15'h1d67: char_row_bitmap <= 16'b0000000000000000;
		15'h1d68: char_row_bitmap <= 16'b0000000000000000;
		15'h1d69: char_row_bitmap <= 16'b0000000000000000;
		15'h1d6a: char_row_bitmap <= 16'b0000000000000000;
		15'h1d6b: char_row_bitmap <= 16'b0000000000000000;
		15'h1d6c: char_row_bitmap <= 16'b0000000000000000;
		15'h1d6d: char_row_bitmap <= 16'b0000000000000000;
		15'h1d6e: char_row_bitmap <= 16'b0000000000000000;
		15'h1d6f: char_row_bitmap <= 16'b0000000000000000;
		15'h1d70: char_row_bitmap <= 16'b0000000000000000;
		15'h1d71: char_row_bitmap <= 16'b0000000000000000;
		15'h1d72: char_row_bitmap <= 16'b0000000000000000;
		15'h1d73: char_row_bitmap <= 16'b0000000000000000;
		15'h1d74: char_row_bitmap <= 16'b0000000000000000;
		15'h1d75: char_row_bitmap <= 16'b0000000000000000;
		15'h1d76: char_row_bitmap <= 16'b0000000000000000;
		15'h1d77: char_row_bitmap <= 16'b0000000000000000;
		15'h1d78: char_row_bitmap <= 16'b0000000000000000;
		15'h1d79: char_row_bitmap <= 16'b0000000000000000;
		15'h1d7a: char_row_bitmap <= 16'b0000000000000000;
		15'h1d7b: char_row_bitmap <= 16'b0000000000000000;
		15'h1d7c: char_row_bitmap <= 16'b0000000000000000;
		15'h1d7d: char_row_bitmap <= 16'b0000000000000000;
		15'h1d7e: char_row_bitmap <= 16'b0000000000000000;
		15'h1d7f: char_row_bitmap <= 16'b0000000000000000;
		15'h1d80: char_row_bitmap <= 16'b0000000000000000;
		15'h1d81: char_row_bitmap <= 16'b0000000000000000;
		15'h1d82: char_row_bitmap <= 16'b0000000000000000;
		15'h1d83: char_row_bitmap <= 16'b0000000000000000;
		15'h1d84: char_row_bitmap <= 16'b0000000000000000;
		15'h1d85: char_row_bitmap <= 16'b0000000000000000;
		15'h1d86: char_row_bitmap <= 16'b0000000000000000;
		15'h1d87: char_row_bitmap <= 16'b0000000000000000;
		15'h1d88: char_row_bitmap <= 16'b0000000000000000;
		15'h1d89: char_row_bitmap <= 16'b0000000000000000;
		15'h1d8a: char_row_bitmap <= 16'b0000000000000000;
		15'h1d8b: char_row_bitmap <= 16'b0000000000000000;
		15'h1d8c: char_row_bitmap <= 16'b0000000000000000;
		15'h1d8d: char_row_bitmap <= 16'b0000000000000000;
		15'h1d8e: char_row_bitmap <= 16'b0000000000000000;
		15'h1d8f: char_row_bitmap <= 16'b0000000000000000;
		15'h1d90: char_row_bitmap <= 16'b0000000000000000;
		15'h1d91: char_row_bitmap <= 16'b0000000000000000;
		15'h1d92: char_row_bitmap <= 16'b0000000000000000;
		15'h1d93: char_row_bitmap <= 16'b0000000000000000;
		15'h1d94: char_row_bitmap <= 16'b0000000000000000;
		15'h1d95: char_row_bitmap <= 16'b0000000000000000;
		15'h1d96: char_row_bitmap <= 16'b0000000000000000;
		15'h1d97: char_row_bitmap <= 16'b0000000000000000;
		15'h1d98: char_row_bitmap <= 16'b0000000000000000;
		15'h1d99: char_row_bitmap <= 16'b0000000000000000;
		15'h1d9a: char_row_bitmap <= 16'b0000000000000000;
		15'h1d9b: char_row_bitmap <= 16'b0000000000000000;
		15'h1d9c: char_row_bitmap <= 16'b0000000000000000;
		15'h1d9d: char_row_bitmap <= 16'b0000000000000000;
		15'h1d9e: char_row_bitmap <= 16'b0000000000000000;
		15'h1d9f: char_row_bitmap <= 16'b0000000000000000;
		15'h1da0: char_row_bitmap <= 16'b0000000000000000;
		15'h1da1: char_row_bitmap <= 16'b0000000000000000;
		15'h1da2: char_row_bitmap <= 16'b0000000000000000;
		15'h1da3: char_row_bitmap <= 16'b0000000000000000;
		15'h1da4: char_row_bitmap <= 16'b0000000000000000;
		15'h1da5: char_row_bitmap <= 16'b0000000000000000;
		15'h1da6: char_row_bitmap <= 16'b0000000000000000;
		15'h1da7: char_row_bitmap <= 16'b0000000000000000;
		15'h1da8: char_row_bitmap <= 16'b0000000000000000;
		15'h1da9: char_row_bitmap <= 16'b0000000000000000;
		15'h1daa: char_row_bitmap <= 16'b0000000000000000;
		15'h1dab: char_row_bitmap <= 16'b0000000000000000;
		15'h1dac: char_row_bitmap <= 16'b0000000000000000;
		15'h1dad: char_row_bitmap <= 16'b0000000000000000;
		15'h1dae: char_row_bitmap <= 16'b0000000000000000;
		15'h1daf: char_row_bitmap <= 16'b0000000000000000;
		15'h1db0: char_row_bitmap <= 16'b0000000000000000;
		15'h1db1: char_row_bitmap <= 16'b0000000000000000;
		15'h1db2: char_row_bitmap <= 16'b0000000000000000;
		15'h1db3: char_row_bitmap <= 16'b0000000000000000;
		15'h1db4: char_row_bitmap <= 16'b0000000000000000;
		15'h1db5: char_row_bitmap <= 16'b0000000000000000;
		15'h1db6: char_row_bitmap <= 16'b0000000000000000;
		15'h1db7: char_row_bitmap <= 16'b0000000000000000;
		15'h1db8: char_row_bitmap <= 16'b0000000000000000;
		15'h1db9: char_row_bitmap <= 16'b0000000000000000;
		15'h1dba: char_row_bitmap <= 16'b0000000000000000;
		15'h1dbb: char_row_bitmap <= 16'b0000000000000000;
		15'h1dbc: char_row_bitmap <= 16'b0000000000000000;
		15'h1dbd: char_row_bitmap <= 16'b0000000000000000;
		15'h1dbe: char_row_bitmap <= 16'b0000000000000000;
		15'h1dbf: char_row_bitmap <= 16'b0000000000000000;
		15'h1dc0: char_row_bitmap <= 16'b0000000000000000;
		15'h1dc1: char_row_bitmap <= 16'b0000000000000000;
		15'h1dc2: char_row_bitmap <= 16'b0000000000000000;
		15'h1dc3: char_row_bitmap <= 16'b0000000000000000;
		15'h1dc4: char_row_bitmap <= 16'b0000000000000000;
		15'h1dc5: char_row_bitmap <= 16'b0000000000000000;
		15'h1dc6: char_row_bitmap <= 16'b0000000000000000;
		15'h1dc7: char_row_bitmap <= 16'b0000000000000000;
		15'h1dc8: char_row_bitmap <= 16'b0000000000000000;
		15'h1dc9: char_row_bitmap <= 16'b0000000000000000;
		15'h1dca: char_row_bitmap <= 16'b0000000000000000;
		15'h1dcb: char_row_bitmap <= 16'b0000000000000000;
		15'h1dcc: char_row_bitmap <= 16'b0000000000000000;
		15'h1dcd: char_row_bitmap <= 16'b0000000000000000;
		15'h1dce: char_row_bitmap <= 16'b0000000000000000;
		15'h1dcf: char_row_bitmap <= 16'b0000000000000000;
		15'h1dd0: char_row_bitmap <= 16'b0000000000000000;
		15'h1dd1: char_row_bitmap <= 16'b0000000000000000;
		15'h1dd2: char_row_bitmap <= 16'b0000000000000000;
		15'h1dd3: char_row_bitmap <= 16'b0000000000000000;
		15'h1dd4: char_row_bitmap <= 16'b0000000000000000;
		15'h1dd5: char_row_bitmap <= 16'b0000000000000000;
		15'h1dd6: char_row_bitmap <= 16'b0000000000000000;
		15'h1dd7: char_row_bitmap <= 16'b0000000000000000;
		15'h1dd8: char_row_bitmap <= 16'b0000000000000000;
		15'h1dd9: char_row_bitmap <= 16'b0000000000000000;
		15'h1dda: char_row_bitmap <= 16'b0000000000000000;
		15'h1ddb: char_row_bitmap <= 16'b0000000000000000;
		15'h1ddc: char_row_bitmap <= 16'b0000000000000000;
		15'h1ddd: char_row_bitmap <= 16'b0000000000000000;
		15'h1dde: char_row_bitmap <= 16'b0000000000000000;
		15'h1ddf: char_row_bitmap <= 16'b0000000000000000;
		15'h1de0: char_row_bitmap <= 16'b0000000000000000;
		15'h1de1: char_row_bitmap <= 16'b0000000000000000;
		15'h1de2: char_row_bitmap <= 16'b0000000000000000;
		15'h1de3: char_row_bitmap <= 16'b0000000000000000;
		15'h1de4: char_row_bitmap <= 16'b0000000000000000;
		15'h1de5: char_row_bitmap <= 16'b0000000000000000;
		15'h1de6: char_row_bitmap <= 16'b0000000000000000;
		15'h1de7: char_row_bitmap <= 16'b0000000000000000;
		15'h1de8: char_row_bitmap <= 16'b0000000000000000;
		15'h1de9: char_row_bitmap <= 16'b0000000000000000;
		15'h1dea: char_row_bitmap <= 16'b0000000000000000;
		15'h1deb: char_row_bitmap <= 16'b0000000000000000;
		15'h1dec: char_row_bitmap <= 16'b0000000000000000;
		15'h1ded: char_row_bitmap <= 16'b0000000000000000;
		15'h1dee: char_row_bitmap <= 16'b0000000000000000;
		15'h1def: char_row_bitmap <= 16'b0000000000000000;
		15'h1df0: char_row_bitmap <= 16'b0000000000000000;
		15'h1df1: char_row_bitmap <= 16'b0000000000000000;
		15'h1df2: char_row_bitmap <= 16'b0000000000000000;
		15'h1df3: char_row_bitmap <= 16'b0000000000000000;
		15'h1df4: char_row_bitmap <= 16'b0000000000000000;
		15'h1df5: char_row_bitmap <= 16'b0000000000000000;
		15'h1df6: char_row_bitmap <= 16'b0000000000000000;
		15'h1df7: char_row_bitmap <= 16'b0000000000000000;
		15'h1df8: char_row_bitmap <= 16'b0000000000000000;
		15'h1df9: char_row_bitmap <= 16'b0000000000000000;
		15'h1dfa: char_row_bitmap <= 16'b0000000000000000;
		15'h1dfb: char_row_bitmap <= 16'b0000000000000000;
		15'h1dfc: char_row_bitmap <= 16'b0000000000000000;
		15'h1dfd: char_row_bitmap <= 16'b0000000000000000;
		15'h1dfe: char_row_bitmap <= 16'b0000000000000000;
		15'h1dff: char_row_bitmap <= 16'b0000000000000000;
		15'h1e00: char_row_bitmap <= 16'b0000000000000000;
		15'h1e01: char_row_bitmap <= 16'b0000000000000000;
		15'h1e02: char_row_bitmap <= 16'b0000000000000000;
		15'h1e03: char_row_bitmap <= 16'b0000000000000000;
		15'h1e04: char_row_bitmap <= 16'b0000000000000000;
		15'h1e05: char_row_bitmap <= 16'b0000000000000000;
		15'h1e06: char_row_bitmap <= 16'b0000000000000000;
		15'h1e07: char_row_bitmap <= 16'b0000000000000000;
		15'h1e08: char_row_bitmap <= 16'b0000000000000000;
		15'h1e09: char_row_bitmap <= 16'b0000000110000000;
		15'h1e0a: char_row_bitmap <= 16'b0000000110000000;
		15'h1e0b: char_row_bitmap <= 16'b0000000000000000;
		15'h1e0c: char_row_bitmap <= 16'b0000000000000000;
		15'h1e0d: char_row_bitmap <= 16'b0000000000000000;
		15'h1e0e: char_row_bitmap <= 16'b0000000000000000;
		15'h1e0f: char_row_bitmap <= 16'b0000000000000000;
		15'h1e10: char_row_bitmap <= 16'b0000000000000000;
		15'h1e11: char_row_bitmap <= 16'b0000000000000000;
		15'h1e12: char_row_bitmap <= 16'b0000000000000000;
		15'h1e13: char_row_bitmap <= 16'b0000000000000000;
		15'h1e14: char_row_bitmap <= 16'b0000000110000000;
		15'h1e15: char_row_bitmap <= 16'b0000000110000000;
		15'h1e16: char_row_bitmap <= 16'b0000000110000000;
		15'h1e17: char_row_bitmap <= 16'b0000000110000000;
		15'h1e18: char_row_bitmap <= 16'b0000000110000000;
		15'h1e19: char_row_bitmap <= 16'b0000000110000000;
		15'h1e1a: char_row_bitmap <= 16'b0000000110000000;
		15'h1e1b: char_row_bitmap <= 16'b0000000110000000;
		15'h1e1c: char_row_bitmap <= 16'b0000000110000000;
		15'h1e1d: char_row_bitmap <= 16'b0000000110000000;
		15'h1e1e: char_row_bitmap <= 16'b0000000110000000;
		15'h1e1f: char_row_bitmap <= 16'b0000000000000000;
		15'h1e20: char_row_bitmap <= 16'b0000000000000000;
		15'h1e21: char_row_bitmap <= 16'b0000000000000000;
		15'h1e22: char_row_bitmap <= 16'b0000000000000000;
		15'h1e23: char_row_bitmap <= 16'b0000000000000000;
		15'h1e24: char_row_bitmap <= 16'b0000000000000000;
		15'h1e25: char_row_bitmap <= 16'b0000000000000000;
		15'h1e26: char_row_bitmap <= 16'b0000000000000000;
		15'h1e27: char_row_bitmap <= 16'b0000000000000000;
		15'h1e28: char_row_bitmap <= 16'b0000000000000000;
		15'h1e29: char_row_bitmap <= 16'b0000000000000000;
		15'h1e2a: char_row_bitmap <= 16'b0000000000000000;
		15'h1e2b: char_row_bitmap <= 16'b0000000000000000;
		15'h1e2c: char_row_bitmap <= 16'b0000000000000000;
		15'h1e2d: char_row_bitmap <= 16'b0000000000000000;
		15'h1e2e: char_row_bitmap <= 16'b0000000000000000;
		15'h1e2f: char_row_bitmap <= 16'b0000000000000000;
		15'h1e30: char_row_bitmap <= 16'b0000000000000000;
		15'h1e31: char_row_bitmap <= 16'b0000000111111111;
		15'h1e32: char_row_bitmap <= 16'b0000000111111111;
		15'h1e33: char_row_bitmap <= 16'b0000000000000000;
		15'h1e34: char_row_bitmap <= 16'b0000000000000000;
		15'h1e35: char_row_bitmap <= 16'b0000000000000000;
		15'h1e36: char_row_bitmap <= 16'b0000000000000000;
		15'h1e37: char_row_bitmap <= 16'b0000000000000000;
		15'h1e38: char_row_bitmap <= 16'b0000000000000000;
		15'h1e39: char_row_bitmap <= 16'b0000000000000000;
		15'h1e3a: char_row_bitmap <= 16'b0000000000000000;
		15'h1e3b: char_row_bitmap <= 16'b0000000000000000;
		15'h1e3c: char_row_bitmap <= 16'b0000000110000000;
		15'h1e3d: char_row_bitmap <= 16'b0000000110000000;
		15'h1e3e: char_row_bitmap <= 16'b0000000110000000;
		15'h1e3f: char_row_bitmap <= 16'b0000000110000000;
		15'h1e40: char_row_bitmap <= 16'b0000000110000000;
		15'h1e41: char_row_bitmap <= 16'b0000000110000000;
		15'h1e42: char_row_bitmap <= 16'b0000000110000000;
		15'h1e43: char_row_bitmap <= 16'b0000000110000000;
		15'h1e44: char_row_bitmap <= 16'b0000000110000000;
		15'h1e45: char_row_bitmap <= 16'b0000000111111111;
		15'h1e46: char_row_bitmap <= 16'b0000000111111111;
		15'h1e47: char_row_bitmap <= 16'b0000000000000000;
		15'h1e48: char_row_bitmap <= 16'b0000000000000000;
		15'h1e49: char_row_bitmap <= 16'b0000000000000000;
		15'h1e4a: char_row_bitmap <= 16'b0000000000000000;
		15'h1e4b: char_row_bitmap <= 16'b0000000000000000;
		15'h1e4c: char_row_bitmap <= 16'b0000000000000000;
		15'h1e4d: char_row_bitmap <= 16'b0000000000000000;
		15'h1e4e: char_row_bitmap <= 16'b0000000000000000;
		15'h1e4f: char_row_bitmap <= 16'b0000000000000000;
		15'h1e50: char_row_bitmap <= 16'b0000000000000000;
		15'h1e51: char_row_bitmap <= 16'b0000000000000000;
		15'h1e52: char_row_bitmap <= 16'b0000000000000000;
		15'h1e53: char_row_bitmap <= 16'b0000000000000000;
		15'h1e54: char_row_bitmap <= 16'b0000000000000000;
		15'h1e55: char_row_bitmap <= 16'b0000000000000000;
		15'h1e56: char_row_bitmap <= 16'b0000000000000000;
		15'h1e57: char_row_bitmap <= 16'b0000000000000000;
		15'h1e58: char_row_bitmap <= 16'b0000000000000000;
		15'h1e59: char_row_bitmap <= 16'b0000000110000000;
		15'h1e5a: char_row_bitmap <= 16'b0000000110000000;
		15'h1e5b: char_row_bitmap <= 16'b0000000110000000;
		15'h1e5c: char_row_bitmap <= 16'b0000000110000000;
		15'h1e5d: char_row_bitmap <= 16'b0000000110000000;
		15'h1e5e: char_row_bitmap <= 16'b0000000110000000;
		15'h1e5f: char_row_bitmap <= 16'b0000000110000000;
		15'h1e60: char_row_bitmap <= 16'b0000000110000000;
		15'h1e61: char_row_bitmap <= 16'b0000000110000000;
		15'h1e62: char_row_bitmap <= 16'b0000000110000000;
		15'h1e63: char_row_bitmap <= 16'b0000000110000000;
		15'h1e64: char_row_bitmap <= 16'b0000000110000000;
		15'h1e65: char_row_bitmap <= 16'b0000000110000000;
		15'h1e66: char_row_bitmap <= 16'b0000000110000000;
		15'h1e67: char_row_bitmap <= 16'b0000000110000000;
		15'h1e68: char_row_bitmap <= 16'b0000000110000000;
		15'h1e69: char_row_bitmap <= 16'b0000000110000000;
		15'h1e6a: char_row_bitmap <= 16'b0000000110000000;
		15'h1e6b: char_row_bitmap <= 16'b0000000110000000;
		15'h1e6c: char_row_bitmap <= 16'b0000000110000000;
		15'h1e6d: char_row_bitmap <= 16'b0000000110000000;
		15'h1e6e: char_row_bitmap <= 16'b0000000110000000;
		15'h1e6f: char_row_bitmap <= 16'b0000000110000000;
		15'h1e70: char_row_bitmap <= 16'b0000000110000000;
		15'h1e71: char_row_bitmap <= 16'b0000000110000000;
		15'h1e72: char_row_bitmap <= 16'b0000000110000000;
		15'h1e73: char_row_bitmap <= 16'b0000000110000000;
		15'h1e74: char_row_bitmap <= 16'b0000000110000000;
		15'h1e75: char_row_bitmap <= 16'b0000000110000000;
		15'h1e76: char_row_bitmap <= 16'b0000000110000000;
		15'h1e77: char_row_bitmap <= 16'b0000000110000000;
		15'h1e78: char_row_bitmap <= 16'b0000000000000000;
		15'h1e79: char_row_bitmap <= 16'b0000000000000000;
		15'h1e7a: char_row_bitmap <= 16'b0000000000000000;
		15'h1e7b: char_row_bitmap <= 16'b0000000000000000;
		15'h1e7c: char_row_bitmap <= 16'b0000000000000000;
		15'h1e7d: char_row_bitmap <= 16'b0000000000000000;
		15'h1e7e: char_row_bitmap <= 16'b0000000000000000;
		15'h1e7f: char_row_bitmap <= 16'b0000000000000000;
		15'h1e80: char_row_bitmap <= 16'b0000000000000000;
		15'h1e81: char_row_bitmap <= 16'b0000000111111111;
		15'h1e82: char_row_bitmap <= 16'b0000000111111111;
		15'h1e83: char_row_bitmap <= 16'b0000000110000000;
		15'h1e84: char_row_bitmap <= 16'b0000000110000000;
		15'h1e85: char_row_bitmap <= 16'b0000000110000000;
		15'h1e86: char_row_bitmap <= 16'b0000000110000000;
		15'h1e87: char_row_bitmap <= 16'b0000000110000000;
		15'h1e88: char_row_bitmap <= 16'b0000000110000000;
		15'h1e89: char_row_bitmap <= 16'b0000000110000000;
		15'h1e8a: char_row_bitmap <= 16'b0000000110000000;
		15'h1e8b: char_row_bitmap <= 16'b0000000110000000;
		15'h1e8c: char_row_bitmap <= 16'b0000000110000000;
		15'h1e8d: char_row_bitmap <= 16'b0000000110000000;
		15'h1e8e: char_row_bitmap <= 16'b0000000110000000;
		15'h1e8f: char_row_bitmap <= 16'b0000000110000000;
		15'h1e90: char_row_bitmap <= 16'b0000000110000000;
		15'h1e91: char_row_bitmap <= 16'b0000000110000000;
		15'h1e92: char_row_bitmap <= 16'b0000000110000000;
		15'h1e93: char_row_bitmap <= 16'b0000000110000000;
		15'h1e94: char_row_bitmap <= 16'b0000000110000000;
		15'h1e95: char_row_bitmap <= 16'b0000000111111111;
		15'h1e96: char_row_bitmap <= 16'b0000000111111111;
		15'h1e97: char_row_bitmap <= 16'b0000000110000000;
		15'h1e98: char_row_bitmap <= 16'b0000000110000000;
		15'h1e99: char_row_bitmap <= 16'b0000000110000000;
		15'h1e9a: char_row_bitmap <= 16'b0000000110000000;
		15'h1e9b: char_row_bitmap <= 16'b0000000110000000;
		15'h1e9c: char_row_bitmap <= 16'b0000000110000000;
		15'h1e9d: char_row_bitmap <= 16'b0000000110000000;
		15'h1e9e: char_row_bitmap <= 16'b0000000110000000;
		15'h1e9f: char_row_bitmap <= 16'b0000000110000000;
		15'h1ea0: char_row_bitmap <= 16'b0000000000000000;
		15'h1ea1: char_row_bitmap <= 16'b0000000000000000;
		15'h1ea2: char_row_bitmap <= 16'b0000000000000000;
		15'h1ea3: char_row_bitmap <= 16'b0000000000000000;
		15'h1ea4: char_row_bitmap <= 16'b0000000000000000;
		15'h1ea5: char_row_bitmap <= 16'b0000000000000000;
		15'h1ea6: char_row_bitmap <= 16'b0000000000000000;
		15'h1ea7: char_row_bitmap <= 16'b0000000000000000;
		15'h1ea8: char_row_bitmap <= 16'b0000000000000000;
		15'h1ea9: char_row_bitmap <= 16'b1111111110000000;
		15'h1eaa: char_row_bitmap <= 16'b1111111110000000;
		15'h1eab: char_row_bitmap <= 16'b0000000000000000;
		15'h1eac: char_row_bitmap <= 16'b0000000000000000;
		15'h1ead: char_row_bitmap <= 16'b0000000000000000;
		15'h1eae: char_row_bitmap <= 16'b0000000000000000;
		15'h1eaf: char_row_bitmap <= 16'b0000000000000000;
		15'h1eb0: char_row_bitmap <= 16'b0000000000000000;
		15'h1eb1: char_row_bitmap <= 16'b0000000000000000;
		15'h1eb2: char_row_bitmap <= 16'b0000000000000000;
		15'h1eb3: char_row_bitmap <= 16'b0000000000000000;
		15'h1eb4: char_row_bitmap <= 16'b0000000110000000;
		15'h1eb5: char_row_bitmap <= 16'b0000000110000000;
		15'h1eb6: char_row_bitmap <= 16'b0000000110000000;
		15'h1eb7: char_row_bitmap <= 16'b0000000110000000;
		15'h1eb8: char_row_bitmap <= 16'b0000000110000000;
		15'h1eb9: char_row_bitmap <= 16'b0000000110000000;
		15'h1eba: char_row_bitmap <= 16'b0000000110000000;
		15'h1ebb: char_row_bitmap <= 16'b0000000110000000;
		15'h1ebc: char_row_bitmap <= 16'b0000000110000000;
		15'h1ebd: char_row_bitmap <= 16'b1111111110000000;
		15'h1ebe: char_row_bitmap <= 16'b1111111110000000;
		15'h1ebf: char_row_bitmap <= 16'b0000000000000000;
		15'h1ec0: char_row_bitmap <= 16'b0000000000000000;
		15'h1ec1: char_row_bitmap <= 16'b0000000000000000;
		15'h1ec2: char_row_bitmap <= 16'b0000000000000000;
		15'h1ec3: char_row_bitmap <= 16'b0000000000000000;
		15'h1ec4: char_row_bitmap <= 16'b0000000000000000;
		15'h1ec5: char_row_bitmap <= 16'b0000000000000000;
		15'h1ec6: char_row_bitmap <= 16'b0000000000000000;
		15'h1ec7: char_row_bitmap <= 16'b0000000000000000;
		15'h1ec8: char_row_bitmap <= 16'b0000000000000000;
		15'h1ec9: char_row_bitmap <= 16'b0000000000000000;
		15'h1eca: char_row_bitmap <= 16'b0000000000000000;
		15'h1ecb: char_row_bitmap <= 16'b0000000000000000;
		15'h1ecc: char_row_bitmap <= 16'b0000000000000000;
		15'h1ecd: char_row_bitmap <= 16'b0000000000000000;
		15'h1ece: char_row_bitmap <= 16'b0000000000000000;
		15'h1ecf: char_row_bitmap <= 16'b0000000000000000;
		15'h1ed0: char_row_bitmap <= 16'b0000000000000000;
		15'h1ed1: char_row_bitmap <= 16'b1111111111111111;
		15'h1ed2: char_row_bitmap <= 16'b1111111111111111;
		15'h1ed3: char_row_bitmap <= 16'b0000000000000000;
		15'h1ed4: char_row_bitmap <= 16'b0000000000000000;
		15'h1ed5: char_row_bitmap <= 16'b0000000000000000;
		15'h1ed6: char_row_bitmap <= 16'b0000000000000000;
		15'h1ed7: char_row_bitmap <= 16'b0000000000000000;
		15'h1ed8: char_row_bitmap <= 16'b0000000000000000;
		15'h1ed9: char_row_bitmap <= 16'b0000000000000000;
		15'h1eda: char_row_bitmap <= 16'b0000000000000000;
		15'h1edb: char_row_bitmap <= 16'b0000000000000000;
		15'h1edc: char_row_bitmap <= 16'b0000000110000000;
		15'h1edd: char_row_bitmap <= 16'b0000000110000000;
		15'h1ede: char_row_bitmap <= 16'b0000000110000000;
		15'h1edf: char_row_bitmap <= 16'b0000000110000000;
		15'h1ee0: char_row_bitmap <= 16'b0000000110000000;
		15'h1ee1: char_row_bitmap <= 16'b0000000110000000;
		15'h1ee2: char_row_bitmap <= 16'b0000000110000000;
		15'h1ee3: char_row_bitmap <= 16'b0000000110000000;
		15'h1ee4: char_row_bitmap <= 16'b0000000110000000;
		15'h1ee5: char_row_bitmap <= 16'b1111111111111111;
		15'h1ee6: char_row_bitmap <= 16'b1111111111111111;
		15'h1ee7: char_row_bitmap <= 16'b0000000000000000;
		15'h1ee8: char_row_bitmap <= 16'b0000000000000000;
		15'h1ee9: char_row_bitmap <= 16'b0000000000000000;
		15'h1eea: char_row_bitmap <= 16'b0000000000000000;
		15'h1eeb: char_row_bitmap <= 16'b0000000000000000;
		15'h1eec: char_row_bitmap <= 16'b0000000000000000;
		15'h1eed: char_row_bitmap <= 16'b0000000000000000;
		15'h1eee: char_row_bitmap <= 16'b0000000000000000;
		15'h1eef: char_row_bitmap <= 16'b0000000000000000;
		15'h1ef0: char_row_bitmap <= 16'b0000000000000000;
		15'h1ef1: char_row_bitmap <= 16'b0000000000000000;
		15'h1ef2: char_row_bitmap <= 16'b0000000000000000;
		15'h1ef3: char_row_bitmap <= 16'b0000000000000000;
		15'h1ef4: char_row_bitmap <= 16'b0000000000000000;
		15'h1ef5: char_row_bitmap <= 16'b0000000000000000;
		15'h1ef6: char_row_bitmap <= 16'b0000000000000000;
		15'h1ef7: char_row_bitmap <= 16'b0000000000000000;
		15'h1ef8: char_row_bitmap <= 16'b0000000000000000;
		15'h1ef9: char_row_bitmap <= 16'b1111111110000000;
		15'h1efa: char_row_bitmap <= 16'b1111111110000000;
		15'h1efb: char_row_bitmap <= 16'b0000000110000000;
		15'h1efc: char_row_bitmap <= 16'b0000000110000000;
		15'h1efd: char_row_bitmap <= 16'b0000000110000000;
		15'h1efe: char_row_bitmap <= 16'b0000000110000000;
		15'h1eff: char_row_bitmap <= 16'b0000000110000000;
		15'h1f00: char_row_bitmap <= 16'b0000000110000000;
		15'h1f01: char_row_bitmap <= 16'b0000000110000000;
		15'h1f02: char_row_bitmap <= 16'b0000000110000000;
		15'h1f03: char_row_bitmap <= 16'b0000000110000000;
		15'h1f04: char_row_bitmap <= 16'b0000000110000000;
		15'h1f05: char_row_bitmap <= 16'b0000000110000000;
		15'h1f06: char_row_bitmap <= 16'b0000000110000000;
		15'h1f07: char_row_bitmap <= 16'b0000000110000000;
		15'h1f08: char_row_bitmap <= 16'b0000000110000000;
		15'h1f09: char_row_bitmap <= 16'b0000000110000000;
		15'h1f0a: char_row_bitmap <= 16'b0000000110000000;
		15'h1f0b: char_row_bitmap <= 16'b0000000110000000;
		15'h1f0c: char_row_bitmap <= 16'b0000000110000000;
		15'h1f0d: char_row_bitmap <= 16'b1111111110000000;
		15'h1f0e: char_row_bitmap <= 16'b1111111110000000;
		15'h1f0f: char_row_bitmap <= 16'b0000000110000000;
		15'h1f10: char_row_bitmap <= 16'b0000000110000000;
		15'h1f11: char_row_bitmap <= 16'b0000000110000000;
		15'h1f12: char_row_bitmap <= 16'b0000000110000000;
		15'h1f13: char_row_bitmap <= 16'b0000000110000000;
		15'h1f14: char_row_bitmap <= 16'b0000000110000000;
		15'h1f15: char_row_bitmap <= 16'b0000000110000000;
		15'h1f16: char_row_bitmap <= 16'b0000000110000000;
		15'h1f17: char_row_bitmap <= 16'b0000000110000000;
		15'h1f18: char_row_bitmap <= 16'b0000000000000000;
		15'h1f19: char_row_bitmap <= 16'b0000000000000000;
		15'h1f1a: char_row_bitmap <= 16'b0000000000000000;
		15'h1f1b: char_row_bitmap <= 16'b0000000000000000;
		15'h1f1c: char_row_bitmap <= 16'b0000000000000000;
		15'h1f1d: char_row_bitmap <= 16'b0000000000000000;
		15'h1f1e: char_row_bitmap <= 16'b0000000000000000;
		15'h1f1f: char_row_bitmap <= 16'b0000000000000000;
		15'h1f20: char_row_bitmap <= 16'b0000000000000000;
		15'h1f21: char_row_bitmap <= 16'b1111111111111111;
		15'h1f22: char_row_bitmap <= 16'b1111111111111111;
		15'h1f23: char_row_bitmap <= 16'b0000000110000000;
		15'h1f24: char_row_bitmap <= 16'b0000000110000000;
		15'h1f25: char_row_bitmap <= 16'b0000000110000000;
		15'h1f26: char_row_bitmap <= 16'b0000000110000000;
		15'h1f27: char_row_bitmap <= 16'b0000000110000000;
		15'h1f28: char_row_bitmap <= 16'b0000000110000000;
		15'h1f29: char_row_bitmap <= 16'b0000000110000000;
		15'h1f2a: char_row_bitmap <= 16'b0000000110000000;
		15'h1f2b: char_row_bitmap <= 16'b0000000110000000;
		15'h1f2c: char_row_bitmap <= 16'b0000000110000000;
		15'h1f2d: char_row_bitmap <= 16'b0000000110000000;
		15'h1f2e: char_row_bitmap <= 16'b0000000110000000;
		15'h1f2f: char_row_bitmap <= 16'b0000000110000000;
		15'h1f30: char_row_bitmap <= 16'b0000000110000000;
		15'h1f31: char_row_bitmap <= 16'b0000000110000000;
		15'h1f32: char_row_bitmap <= 16'b0000000110000000;
		15'h1f33: char_row_bitmap <= 16'b0000000110000000;
		15'h1f34: char_row_bitmap <= 16'b0000000110000000;
		15'h1f35: char_row_bitmap <= 16'b1111111111111111;
		15'h1f36: char_row_bitmap <= 16'b1111111111111111;
		15'h1f37: char_row_bitmap <= 16'b0000000110000000;
		15'h1f38: char_row_bitmap <= 16'b0000000110000000;
		15'h1f39: char_row_bitmap <= 16'b0000000110000000;
		15'h1f3a: char_row_bitmap <= 16'b0000000110000000;
		15'h1f3b: char_row_bitmap <= 16'b0000000110000000;
		15'h1f3c: char_row_bitmap <= 16'b0000000110000000;
		15'h1f3d: char_row_bitmap <= 16'b0000000110000000;
		15'h1f3e: char_row_bitmap <= 16'b0000000110000000;
		15'h1f3f: char_row_bitmap <= 16'b0000000110000000;
		15'h1f40: char_row_bitmap <= 16'b0000000000000000;
		15'h1f41: char_row_bitmap <= 16'b0000000000000000;
		15'h1f42: char_row_bitmap <= 16'b0000000000000000;
		15'h1f43: char_row_bitmap <= 16'b0000000000000000;
		15'h1f44: char_row_bitmap <= 16'b0000000000000000;
		15'h1f45: char_row_bitmap <= 16'b0000000000000000;
		15'h1f46: char_row_bitmap <= 16'b0000000000000000;
		15'h1f47: char_row_bitmap <= 16'b0000000000000000;
		15'h1f48: char_row_bitmap <= 16'b0000001111000000;
		15'h1f49: char_row_bitmap <= 16'b0000001001000000;
		15'h1f4a: char_row_bitmap <= 16'b0000001001000000;
		15'h1f4b: char_row_bitmap <= 16'b0000001111000000;
		15'h1f4c: char_row_bitmap <= 16'b0000000000000000;
		15'h1f4d: char_row_bitmap <= 16'b0000000000000000;
		15'h1f4e: char_row_bitmap <= 16'b0000000000000000;
		15'h1f4f: char_row_bitmap <= 16'b0000000000000000;
		15'h1f50: char_row_bitmap <= 16'b0000000000000000;
		15'h1f51: char_row_bitmap <= 16'b0000000000000000;
		15'h1f52: char_row_bitmap <= 16'b0000000000000000;
		15'h1f53: char_row_bitmap <= 16'b0000000000000000;
		15'h1f54: char_row_bitmap <= 16'b0000001001000000;
		15'h1f55: char_row_bitmap <= 16'b0000001001000000;
		15'h1f56: char_row_bitmap <= 16'b0000001001000000;
		15'h1f57: char_row_bitmap <= 16'b0000001001000000;
		15'h1f58: char_row_bitmap <= 16'b0000001001000000;
		15'h1f59: char_row_bitmap <= 16'b0000001001000000;
		15'h1f5a: char_row_bitmap <= 16'b0000001001000000;
		15'h1f5b: char_row_bitmap <= 16'b0000001001000000;
		15'h1f5c: char_row_bitmap <= 16'b0000001001000000;
		15'h1f5d: char_row_bitmap <= 16'b0000001001000000;
		15'h1f5e: char_row_bitmap <= 16'b0000001001000000;
		15'h1f5f: char_row_bitmap <= 16'b0000001111000000;
		15'h1f60: char_row_bitmap <= 16'b0000000000000000;
		15'h1f61: char_row_bitmap <= 16'b0000000000000000;
		15'h1f62: char_row_bitmap <= 16'b0000000000000000;
		15'h1f63: char_row_bitmap <= 16'b0000000000000000;
		15'h1f64: char_row_bitmap <= 16'b0000000000000000;
		15'h1f65: char_row_bitmap <= 16'b0000000000000000;
		15'h1f66: char_row_bitmap <= 16'b0000000000000000;
		15'h1f67: char_row_bitmap <= 16'b0000000000000000;
		15'h1f68: char_row_bitmap <= 16'b0000000000000000;
		15'h1f69: char_row_bitmap <= 16'b0000000000000000;
		15'h1f6a: char_row_bitmap <= 16'b0000000000000000;
		15'h1f6b: char_row_bitmap <= 16'b0000000000000000;
		15'h1f6c: char_row_bitmap <= 16'b0000000000000000;
		15'h1f6d: char_row_bitmap <= 16'b0000000000000000;
		15'h1f6e: char_row_bitmap <= 16'b0000000000000000;
		15'h1f6f: char_row_bitmap <= 16'b0000000000000000;
		15'h1f70: char_row_bitmap <= 16'b0000001111111111;
		15'h1f71: char_row_bitmap <= 16'b0000001000000000;
		15'h1f72: char_row_bitmap <= 16'b0000001000000000;
		15'h1f73: char_row_bitmap <= 16'b0000001111111111;
		15'h1f74: char_row_bitmap <= 16'b0000000000000000;
		15'h1f75: char_row_bitmap <= 16'b0000000000000000;
		15'h1f76: char_row_bitmap <= 16'b0000000000000000;
		15'h1f77: char_row_bitmap <= 16'b0000000000000000;
		15'h1f78: char_row_bitmap <= 16'b0000000000000000;
		15'h1f79: char_row_bitmap <= 16'b0000000000000000;
		15'h1f7a: char_row_bitmap <= 16'b0000000000000000;
		15'h1f7b: char_row_bitmap <= 16'b0000000000000000;
		15'h1f7c: char_row_bitmap <= 16'b0000001001000000;
		15'h1f7d: char_row_bitmap <= 16'b0000001001000000;
		15'h1f7e: char_row_bitmap <= 16'b0000001001000000;
		15'h1f7f: char_row_bitmap <= 16'b0000001001000000;
		15'h1f80: char_row_bitmap <= 16'b0000001001000000;
		15'h1f81: char_row_bitmap <= 16'b0000001001000000;
		15'h1f82: char_row_bitmap <= 16'b0000001001000000;
		15'h1f83: char_row_bitmap <= 16'b0000001001000000;
		15'h1f84: char_row_bitmap <= 16'b0000001001111111;
		15'h1f85: char_row_bitmap <= 16'b0000001000000000;
		15'h1f86: char_row_bitmap <= 16'b0000001000000000;
		15'h1f87: char_row_bitmap <= 16'b0000001111111111;
		15'h1f88: char_row_bitmap <= 16'b0000000000000000;
		15'h1f89: char_row_bitmap <= 16'b0000000000000000;
		15'h1f8a: char_row_bitmap <= 16'b0000000000000000;
		15'h1f8b: char_row_bitmap <= 16'b0000000000000000;
		15'h1f8c: char_row_bitmap <= 16'b0000000000000000;
		15'h1f8d: char_row_bitmap <= 16'b0000000000000000;
		15'h1f8e: char_row_bitmap <= 16'b0000000000000000;
		15'h1f8f: char_row_bitmap <= 16'b0000000000000000;
		15'h1f90: char_row_bitmap <= 16'b0000000000000000;
		15'h1f91: char_row_bitmap <= 16'b0000000000000000;
		15'h1f92: char_row_bitmap <= 16'b0000000000000000;
		15'h1f93: char_row_bitmap <= 16'b0000000000000000;
		15'h1f94: char_row_bitmap <= 16'b0000000000000000;
		15'h1f95: char_row_bitmap <= 16'b0000000000000000;
		15'h1f96: char_row_bitmap <= 16'b0000000000000000;
		15'h1f97: char_row_bitmap <= 16'b0000000000000000;
		15'h1f98: char_row_bitmap <= 16'b0000001001000000;
		15'h1f99: char_row_bitmap <= 16'b0000001001000000;
		15'h1f9a: char_row_bitmap <= 16'b0000001001000000;
		15'h1f9b: char_row_bitmap <= 16'b0000001001000000;
		15'h1f9c: char_row_bitmap <= 16'b0000001001000000;
		15'h1f9d: char_row_bitmap <= 16'b0000001001000000;
		15'h1f9e: char_row_bitmap <= 16'b0000001001000000;
		15'h1f9f: char_row_bitmap <= 16'b0000001001000000;
		15'h1fa0: char_row_bitmap <= 16'b0000001001000000;
		15'h1fa1: char_row_bitmap <= 16'b0000001001000000;
		15'h1fa2: char_row_bitmap <= 16'b0000001001000000;
		15'h1fa3: char_row_bitmap <= 16'b0000001001000000;
		15'h1fa4: char_row_bitmap <= 16'b0000001001000000;
		15'h1fa5: char_row_bitmap <= 16'b0000001001000000;
		15'h1fa6: char_row_bitmap <= 16'b0000001001000000;
		15'h1fa7: char_row_bitmap <= 16'b0000001001000000;
		15'h1fa8: char_row_bitmap <= 16'b0000001001000000;
		15'h1fa9: char_row_bitmap <= 16'b0000001001000000;
		15'h1faa: char_row_bitmap <= 16'b0000001001000000;
		15'h1fab: char_row_bitmap <= 16'b0000001001000000;
		15'h1fac: char_row_bitmap <= 16'b0000001001000000;
		15'h1fad: char_row_bitmap <= 16'b0000001001000000;
		15'h1fae: char_row_bitmap <= 16'b0000001001000000;
		15'h1faf: char_row_bitmap <= 16'b0000001001000000;
		15'h1fb0: char_row_bitmap <= 16'b0000001001000000;
		15'h1fb1: char_row_bitmap <= 16'b0000001001000000;
		15'h1fb2: char_row_bitmap <= 16'b0000001001000000;
		15'h1fb3: char_row_bitmap <= 16'b0000001001000000;
		15'h1fb4: char_row_bitmap <= 16'b0000001001000000;
		15'h1fb5: char_row_bitmap <= 16'b0000001001000000;
		15'h1fb6: char_row_bitmap <= 16'b0000001001000000;
		15'h1fb7: char_row_bitmap <= 16'b0000001001000000;
		15'h1fb8: char_row_bitmap <= 16'b0000000000000000;
		15'h1fb9: char_row_bitmap <= 16'b0000000000000000;
		15'h1fba: char_row_bitmap <= 16'b0000000000000000;
		15'h1fbb: char_row_bitmap <= 16'b0000000000000000;
		15'h1fbc: char_row_bitmap <= 16'b0000000000000000;
		15'h1fbd: char_row_bitmap <= 16'b0000000000000000;
		15'h1fbe: char_row_bitmap <= 16'b0000000000000000;
		15'h1fbf: char_row_bitmap <= 16'b0000000000000000;
		15'h1fc0: char_row_bitmap <= 16'b0000001111111111;
		15'h1fc1: char_row_bitmap <= 16'b0000001000000000;
		15'h1fc2: char_row_bitmap <= 16'b0000001000000000;
		15'h1fc3: char_row_bitmap <= 16'b0000001001111111;
		15'h1fc4: char_row_bitmap <= 16'b0000001001000000;
		15'h1fc5: char_row_bitmap <= 16'b0000001001000000;
		15'h1fc6: char_row_bitmap <= 16'b0000001001000000;
		15'h1fc7: char_row_bitmap <= 16'b0000001001000000;
		15'h1fc8: char_row_bitmap <= 16'b0000001001000000;
		15'h1fc9: char_row_bitmap <= 16'b0000001001000000;
		15'h1fca: char_row_bitmap <= 16'b0000001001000000;
		15'h1fcb: char_row_bitmap <= 16'b0000001001000000;
		15'h1fcc: char_row_bitmap <= 16'b0000001001000000;
		15'h1fcd: char_row_bitmap <= 16'b0000001001000000;
		15'h1fce: char_row_bitmap <= 16'b0000001001000000;
		15'h1fcf: char_row_bitmap <= 16'b0000001001000000;
		15'h1fd0: char_row_bitmap <= 16'b0000001001000000;
		15'h1fd1: char_row_bitmap <= 16'b0000001001000000;
		15'h1fd2: char_row_bitmap <= 16'b0000001001000000;
		15'h1fd3: char_row_bitmap <= 16'b0000001001000000;
		15'h1fd4: char_row_bitmap <= 16'b0000001001111111;
		15'h1fd5: char_row_bitmap <= 16'b0000001000000000;
		15'h1fd6: char_row_bitmap <= 16'b0000001000000000;
		15'h1fd7: char_row_bitmap <= 16'b0000001001111111;
		15'h1fd8: char_row_bitmap <= 16'b0000001001000000;
		15'h1fd9: char_row_bitmap <= 16'b0000001001000000;
		15'h1fda: char_row_bitmap <= 16'b0000001001000000;
		15'h1fdb: char_row_bitmap <= 16'b0000001001000000;
		15'h1fdc: char_row_bitmap <= 16'b0000001001000000;
		15'h1fdd: char_row_bitmap <= 16'b0000001001000000;
		15'h1fde: char_row_bitmap <= 16'b0000001001000000;
		15'h1fdf: char_row_bitmap <= 16'b0000001001000000;
		15'h1fe0: char_row_bitmap <= 16'b0000000000000000;
		15'h1fe1: char_row_bitmap <= 16'b0000000000000000;
		15'h1fe2: char_row_bitmap <= 16'b0000000000000000;
		15'h1fe3: char_row_bitmap <= 16'b0000000000000000;
		15'h1fe4: char_row_bitmap <= 16'b0000000000000000;
		15'h1fe5: char_row_bitmap <= 16'b0000000000000000;
		15'h1fe6: char_row_bitmap <= 16'b0000000000000000;
		15'h1fe7: char_row_bitmap <= 16'b0000000000000000;
		15'h1fe8: char_row_bitmap <= 16'b1111111111000000;
		15'h1fe9: char_row_bitmap <= 16'b0000000001000000;
		15'h1fea: char_row_bitmap <= 16'b0000000001000000;
		15'h1feb: char_row_bitmap <= 16'b1111111111000000;
		15'h1fec: char_row_bitmap <= 16'b0000000000000000;
		15'h1fed: char_row_bitmap <= 16'b0000000000000000;
		15'h1fee: char_row_bitmap <= 16'b0000000000000000;
		15'h1fef: char_row_bitmap <= 16'b0000000000000000;
		15'h1ff0: char_row_bitmap <= 16'b0000000000000000;
		15'h1ff1: char_row_bitmap <= 16'b0000000000000000;
		15'h1ff2: char_row_bitmap <= 16'b0000000000000000;
		15'h1ff3: char_row_bitmap <= 16'b0000000000000000;
		15'h1ff4: char_row_bitmap <= 16'b0000001001000000;
		15'h1ff5: char_row_bitmap <= 16'b0000001001000000;
		15'h1ff6: char_row_bitmap <= 16'b0000001001000000;
		15'h1ff7: char_row_bitmap <= 16'b0000001001000000;
		15'h1ff8: char_row_bitmap <= 16'b0000001001000000;
		15'h1ff9: char_row_bitmap <= 16'b0000001001000000;
		15'h1ffa: char_row_bitmap <= 16'b0000001001000000;
		15'h1ffb: char_row_bitmap <= 16'b0000001001000000;
		15'h1ffc: char_row_bitmap <= 16'b1111111001000000;
		15'h1ffd: char_row_bitmap <= 16'b0000000001000000;
		15'h1ffe: char_row_bitmap <= 16'b0000000001000000;
		15'h1fff: char_row_bitmap <= 16'b1111111111000000;
		15'h2000: char_row_bitmap <= 16'b0000000000000000;
		15'h2001: char_row_bitmap <= 16'b0000000000000000;
		15'h2002: char_row_bitmap <= 16'b0000000000000000;
		15'h2003: char_row_bitmap <= 16'b0000000000000000;
		15'h2004: char_row_bitmap <= 16'b0000000000000000;
		15'h2005: char_row_bitmap <= 16'b0000000000000000;
		15'h2006: char_row_bitmap <= 16'b0000000000000000;
		15'h2007: char_row_bitmap <= 16'b0000000000000000;
		15'h2008: char_row_bitmap <= 16'b0000000000000000;
		15'h2009: char_row_bitmap <= 16'b0000000000000000;
		15'h200a: char_row_bitmap <= 16'b0000000000000000;
		15'h200b: char_row_bitmap <= 16'b0000000000000000;
		15'h200c: char_row_bitmap <= 16'b0000000000000000;
		15'h200d: char_row_bitmap <= 16'b0000000000000000;
		15'h200e: char_row_bitmap <= 16'b0000000000000000;
		15'h200f: char_row_bitmap <= 16'b0000000000000000;
		15'h2010: char_row_bitmap <= 16'b1111111111111111;
		15'h2011: char_row_bitmap <= 16'b0000000000000000;
		15'h2012: char_row_bitmap <= 16'b0000000000000000;
		15'h2013: char_row_bitmap <= 16'b1111111111111111;
		15'h2014: char_row_bitmap <= 16'b0000000000000000;
		15'h2015: char_row_bitmap <= 16'b0000000000000000;
		15'h2016: char_row_bitmap <= 16'b0000000000000000;
		15'h2017: char_row_bitmap <= 16'b0000000000000000;
		15'h2018: char_row_bitmap <= 16'b0000000000000000;
		15'h2019: char_row_bitmap <= 16'b0000000000000000;
		15'h201a: char_row_bitmap <= 16'b0000000000000000;
		15'h201b: char_row_bitmap <= 16'b0000000000000000;
		15'h201c: char_row_bitmap <= 16'b0000001001000000;
		15'h201d: char_row_bitmap <= 16'b0000001001000000;
		15'h201e: char_row_bitmap <= 16'b0000001001000000;
		15'h201f: char_row_bitmap <= 16'b0000001001000000;
		15'h2020: char_row_bitmap <= 16'b0000001001000000;
		15'h2021: char_row_bitmap <= 16'b0000001001000000;
		15'h2022: char_row_bitmap <= 16'b0000001001000000;
		15'h2023: char_row_bitmap <= 16'b0000001001000000;
		15'h2024: char_row_bitmap <= 16'b1111111001111111;
		15'h2025: char_row_bitmap <= 16'b0000000000000000;
		15'h2026: char_row_bitmap <= 16'b0000000000000000;
		15'h2027: char_row_bitmap <= 16'b1111111111111111;
		15'h2028: char_row_bitmap <= 16'b0000000000000000;
		15'h2029: char_row_bitmap <= 16'b0000000000000000;
		15'h202a: char_row_bitmap <= 16'b0000000000000000;
		15'h202b: char_row_bitmap <= 16'b0000000000000000;
		15'h202c: char_row_bitmap <= 16'b0000000000000000;
		15'h202d: char_row_bitmap <= 16'b0000000000000000;
		15'h202e: char_row_bitmap <= 16'b0000000000000000;
		15'h202f: char_row_bitmap <= 16'b0000000000000000;
		15'h2030: char_row_bitmap <= 16'b0000000000000000;
		15'h2031: char_row_bitmap <= 16'b0000000000000000;
		15'h2032: char_row_bitmap <= 16'b0000000000000000;
		15'h2033: char_row_bitmap <= 16'b0000000000000000;
		15'h2034: char_row_bitmap <= 16'b0000000000000000;
		15'h2035: char_row_bitmap <= 16'b0000000000000000;
		15'h2036: char_row_bitmap <= 16'b0000000000000000;
		15'h2037: char_row_bitmap <= 16'b0000000000000000;
		15'h2038: char_row_bitmap <= 16'b1111111111000000;
		15'h2039: char_row_bitmap <= 16'b0000000001000000;
		15'h203a: char_row_bitmap <= 16'b0000000001000000;
		15'h203b: char_row_bitmap <= 16'b1111111001000000;
		15'h203c: char_row_bitmap <= 16'b0000001001000000;
		15'h203d: char_row_bitmap <= 16'b0000001001000000;
		15'h203e: char_row_bitmap <= 16'b0000001001000000;
		15'h203f: char_row_bitmap <= 16'b0000001001000000;
		15'h2040: char_row_bitmap <= 16'b0000001001000000;
		15'h2041: char_row_bitmap <= 16'b0000001001000000;
		15'h2042: char_row_bitmap <= 16'b0000001001000000;
		15'h2043: char_row_bitmap <= 16'b0000001001000000;
		15'h2044: char_row_bitmap <= 16'b0000001001000000;
		15'h2045: char_row_bitmap <= 16'b0000001001000000;
		15'h2046: char_row_bitmap <= 16'b0000001001000000;
		15'h2047: char_row_bitmap <= 16'b0000001001000000;
		15'h2048: char_row_bitmap <= 16'b0000001001000000;
		15'h2049: char_row_bitmap <= 16'b0000001001000000;
		15'h204a: char_row_bitmap <= 16'b0000001001000000;
		15'h204b: char_row_bitmap <= 16'b0000001001000000;
		15'h204c: char_row_bitmap <= 16'b1111111001000000;
		15'h204d: char_row_bitmap <= 16'b0000000001000000;
		15'h204e: char_row_bitmap <= 16'b0000000001000000;
		15'h204f: char_row_bitmap <= 16'b1111111001000000;
		15'h2050: char_row_bitmap <= 16'b0000001001000000;
		15'h2051: char_row_bitmap <= 16'b0000001001000000;
		15'h2052: char_row_bitmap <= 16'b0000001001000000;
		15'h2053: char_row_bitmap <= 16'b0000001001000000;
		15'h2054: char_row_bitmap <= 16'b0000001001000000;
		15'h2055: char_row_bitmap <= 16'b0000001001000000;
		15'h2056: char_row_bitmap <= 16'b0000001001000000;
		15'h2057: char_row_bitmap <= 16'b0000001001000000;
		15'h2058: char_row_bitmap <= 16'b0000000000000000;
		15'h2059: char_row_bitmap <= 16'b0000000000000000;
		15'h205a: char_row_bitmap <= 16'b0000000000000000;
		15'h205b: char_row_bitmap <= 16'b0000000000000000;
		15'h205c: char_row_bitmap <= 16'b0000000000000000;
		15'h205d: char_row_bitmap <= 16'b0000000000000000;
		15'h205e: char_row_bitmap <= 16'b0000000000000000;
		15'h205f: char_row_bitmap <= 16'b0000000000000000;
		15'h2060: char_row_bitmap <= 16'b1111111111111111;
		15'h2061: char_row_bitmap <= 16'b0000000000000000;
		15'h2062: char_row_bitmap <= 16'b0000000000000000;
		15'h2063: char_row_bitmap <= 16'b1111111001111111;
		15'h2064: char_row_bitmap <= 16'b0000001001000000;
		15'h2065: char_row_bitmap <= 16'b0000001001000000;
		15'h2066: char_row_bitmap <= 16'b0000001001000000;
		15'h2067: char_row_bitmap <= 16'b0000001001000000;
		15'h2068: char_row_bitmap <= 16'b0000001001000000;
		15'h2069: char_row_bitmap <= 16'b0000001001000000;
		15'h206a: char_row_bitmap <= 16'b0000001001000000;
		15'h206b: char_row_bitmap <= 16'b0000001001000000;
		15'h206c: char_row_bitmap <= 16'b0000001001000000;
		15'h206d: char_row_bitmap <= 16'b0000001001000000;
		15'h206e: char_row_bitmap <= 16'b0000001001000000;
		15'h206f: char_row_bitmap <= 16'b0000001001000000;
		15'h2070: char_row_bitmap <= 16'b0000001001000000;
		15'h2071: char_row_bitmap <= 16'b0000001001000000;
		15'h2072: char_row_bitmap <= 16'b0000001001000000;
		15'h2073: char_row_bitmap <= 16'b0000001001000000;
		15'h2074: char_row_bitmap <= 16'b1111111001111111;
		15'h2075: char_row_bitmap <= 16'b0000000000000000;
		15'h2076: char_row_bitmap <= 16'b0000000000000000;
		15'h2077: char_row_bitmap <= 16'b1111111001111111;
		15'h2078: char_row_bitmap <= 16'b0000001001000000;
		15'h2079: char_row_bitmap <= 16'b0000001001000000;
		15'h207a: char_row_bitmap <= 16'b0000001001000000;
		15'h207b: char_row_bitmap <= 16'b0000001001000000;
		15'h207c: char_row_bitmap <= 16'b0000001001000000;
		15'h207d: char_row_bitmap <= 16'b0000001001000000;
		15'h207e: char_row_bitmap <= 16'b0000001001000000;
		15'h207f: char_row_bitmap <= 16'b0000001001000000;
		15'h2080: char_row_bitmap <= 16'b0000000000000000;
		15'h2081: char_row_bitmap <= 16'b0000000000000000;
		15'h2082: char_row_bitmap <= 16'b0000000000000000;
		15'h2083: char_row_bitmap <= 16'b0000000000000000;
		15'h2084: char_row_bitmap <= 16'b0000000000000000;
		15'h2085: char_row_bitmap <= 16'b0000000000000000;
		15'h2086: char_row_bitmap <= 16'b0000000000000000;
		15'h2087: char_row_bitmap <= 16'b0000000000000000;
		15'h2088: char_row_bitmap <= 16'b0000001111000000;
		15'h2089: char_row_bitmap <= 16'b0000001111000000;
		15'h208a: char_row_bitmap <= 16'b0000001111000000;
		15'h208b: char_row_bitmap <= 16'b0000001111000000;
		15'h208c: char_row_bitmap <= 16'b0000000000000000;
		15'h208d: char_row_bitmap <= 16'b0000000000000000;
		15'h208e: char_row_bitmap <= 16'b0000000000000000;
		15'h208f: char_row_bitmap <= 16'b0000000000000000;
		15'h2090: char_row_bitmap <= 16'b0000000000000000;
		15'h2091: char_row_bitmap <= 16'b0000000000000000;
		15'h2092: char_row_bitmap <= 16'b0000000000000000;
		15'h2093: char_row_bitmap <= 16'b0000000000000000;
		15'h2094: char_row_bitmap <= 16'b0000001111000000;
		15'h2095: char_row_bitmap <= 16'b0000001111000000;
		15'h2096: char_row_bitmap <= 16'b0000001111000000;
		15'h2097: char_row_bitmap <= 16'b0000001111000000;
		15'h2098: char_row_bitmap <= 16'b0000001111000000;
		15'h2099: char_row_bitmap <= 16'b0000001111000000;
		15'h209a: char_row_bitmap <= 16'b0000001111000000;
		15'h209b: char_row_bitmap <= 16'b0000001111000000;
		15'h209c: char_row_bitmap <= 16'b0000001111000000;
		15'h209d: char_row_bitmap <= 16'b0000001111000000;
		15'h209e: char_row_bitmap <= 16'b0000001111000000;
		15'h209f: char_row_bitmap <= 16'b0000001111000000;
		15'h20a0: char_row_bitmap <= 16'b0000000000000000;
		15'h20a1: char_row_bitmap <= 16'b0000000000000000;
		15'h20a2: char_row_bitmap <= 16'b0000000000000000;
		15'h20a3: char_row_bitmap <= 16'b0000000000000000;
		15'h20a4: char_row_bitmap <= 16'b0000000000000000;
		15'h20a5: char_row_bitmap <= 16'b0000000000000000;
		15'h20a6: char_row_bitmap <= 16'b0000000000000000;
		15'h20a7: char_row_bitmap <= 16'b0000000000000000;
		15'h20a8: char_row_bitmap <= 16'b0000000000000000;
		15'h20a9: char_row_bitmap <= 16'b0000000000000000;
		15'h20aa: char_row_bitmap <= 16'b0000000000000000;
		15'h20ab: char_row_bitmap <= 16'b0000000000000000;
		15'h20ac: char_row_bitmap <= 16'b0000000000000000;
		15'h20ad: char_row_bitmap <= 16'b0000000000000000;
		15'h20ae: char_row_bitmap <= 16'b0000000000000000;
		15'h20af: char_row_bitmap <= 16'b0000000000000000;
		15'h20b0: char_row_bitmap <= 16'b0000001111111111;
		15'h20b1: char_row_bitmap <= 16'b0000001111111111;
		15'h20b2: char_row_bitmap <= 16'b0000001111111111;
		15'h20b3: char_row_bitmap <= 16'b0000001111111111;
		15'h20b4: char_row_bitmap <= 16'b0000000000000000;
		15'h20b5: char_row_bitmap <= 16'b0000000000000000;
		15'h20b6: char_row_bitmap <= 16'b0000000000000000;
		15'h20b7: char_row_bitmap <= 16'b0000000000000000;
		15'h20b8: char_row_bitmap <= 16'b0000000000000000;
		15'h20b9: char_row_bitmap <= 16'b0000000000000000;
		15'h20ba: char_row_bitmap <= 16'b0000000000000000;
		15'h20bb: char_row_bitmap <= 16'b0000000000000000;
		15'h20bc: char_row_bitmap <= 16'b0000001111000000;
		15'h20bd: char_row_bitmap <= 16'b0000001111000000;
		15'h20be: char_row_bitmap <= 16'b0000001111000000;
		15'h20bf: char_row_bitmap <= 16'b0000001111000000;
		15'h20c0: char_row_bitmap <= 16'b0000001111000000;
		15'h20c1: char_row_bitmap <= 16'b0000001111000000;
		15'h20c2: char_row_bitmap <= 16'b0000001111000000;
		15'h20c3: char_row_bitmap <= 16'b0000001111000000;
		15'h20c4: char_row_bitmap <= 16'b0000001111111111;
		15'h20c5: char_row_bitmap <= 16'b0000001111111111;
		15'h20c6: char_row_bitmap <= 16'b0000001111111111;
		15'h20c7: char_row_bitmap <= 16'b0000001111111111;
		15'h20c8: char_row_bitmap <= 16'b0000000000000000;
		15'h20c9: char_row_bitmap <= 16'b0000000000000000;
		15'h20ca: char_row_bitmap <= 16'b0000000000000000;
		15'h20cb: char_row_bitmap <= 16'b0000000000000000;
		15'h20cc: char_row_bitmap <= 16'b0000000000000000;
		15'h20cd: char_row_bitmap <= 16'b0000000000000000;
		15'h20ce: char_row_bitmap <= 16'b0000000000000000;
		15'h20cf: char_row_bitmap <= 16'b0000000000000000;
		15'h20d0: char_row_bitmap <= 16'b0000000000000000;
		15'h20d1: char_row_bitmap <= 16'b0000000000000000;
		15'h20d2: char_row_bitmap <= 16'b0000000000000000;
		15'h20d3: char_row_bitmap <= 16'b0000000000000000;
		15'h20d4: char_row_bitmap <= 16'b0000000000000000;
		15'h20d5: char_row_bitmap <= 16'b0000000000000000;
		15'h20d6: char_row_bitmap <= 16'b0000000000000000;
		15'h20d7: char_row_bitmap <= 16'b0000000000000000;
		15'h20d8: char_row_bitmap <= 16'b0000001111000000;
		15'h20d9: char_row_bitmap <= 16'b0000001111000000;
		15'h20da: char_row_bitmap <= 16'b0000001111000000;
		15'h20db: char_row_bitmap <= 16'b0000001111000000;
		15'h20dc: char_row_bitmap <= 16'b0000001111000000;
		15'h20dd: char_row_bitmap <= 16'b0000001111000000;
		15'h20de: char_row_bitmap <= 16'b0000001111000000;
		15'h20df: char_row_bitmap <= 16'b0000001111000000;
		15'h20e0: char_row_bitmap <= 16'b0000001111000000;
		15'h20e1: char_row_bitmap <= 16'b0000001111000000;
		15'h20e2: char_row_bitmap <= 16'b0000001111000000;
		15'h20e3: char_row_bitmap <= 16'b0000001111000000;
		15'h20e4: char_row_bitmap <= 16'b0000001111000000;
		15'h20e5: char_row_bitmap <= 16'b0000001111000000;
		15'h20e6: char_row_bitmap <= 16'b0000001111000000;
		15'h20e7: char_row_bitmap <= 16'b0000001111000000;
		15'h20e8: char_row_bitmap <= 16'b0000001111000000;
		15'h20e9: char_row_bitmap <= 16'b0000001111000000;
		15'h20ea: char_row_bitmap <= 16'b0000001111000000;
		15'h20eb: char_row_bitmap <= 16'b0000001111000000;
		15'h20ec: char_row_bitmap <= 16'b0000001111000000;
		15'h20ed: char_row_bitmap <= 16'b0000001111000000;
		15'h20ee: char_row_bitmap <= 16'b0000001111000000;
		15'h20ef: char_row_bitmap <= 16'b0000001111000000;
		15'h20f0: char_row_bitmap <= 16'b0000001111000000;
		15'h20f1: char_row_bitmap <= 16'b0000001111000000;
		15'h20f2: char_row_bitmap <= 16'b0000001111000000;
		15'h20f3: char_row_bitmap <= 16'b0000001111000000;
		15'h20f4: char_row_bitmap <= 16'b0000001111000000;
		15'h20f5: char_row_bitmap <= 16'b0000001111000000;
		15'h20f6: char_row_bitmap <= 16'b0000001111000000;
		15'h20f7: char_row_bitmap <= 16'b0000001111000000;
		15'h20f8: char_row_bitmap <= 16'b0000000000000000;
		15'h20f9: char_row_bitmap <= 16'b0000000000000000;
		15'h20fa: char_row_bitmap <= 16'b0000000000000000;
		15'h20fb: char_row_bitmap <= 16'b0000000000000000;
		15'h20fc: char_row_bitmap <= 16'b0000000000000000;
		15'h20fd: char_row_bitmap <= 16'b0000000000000000;
		15'h20fe: char_row_bitmap <= 16'b0000000000000000;
		15'h20ff: char_row_bitmap <= 16'b0000000000000000;
		15'h2100: char_row_bitmap <= 16'b0000001111111111;
		15'h2101: char_row_bitmap <= 16'b0000001111111111;
		15'h2102: char_row_bitmap <= 16'b0000001111111111;
		15'h2103: char_row_bitmap <= 16'b0000001111111111;
		15'h2104: char_row_bitmap <= 16'b0000001111000000;
		15'h2105: char_row_bitmap <= 16'b0000001111000000;
		15'h2106: char_row_bitmap <= 16'b0000001111000000;
		15'h2107: char_row_bitmap <= 16'b0000001111000000;
		15'h2108: char_row_bitmap <= 16'b0000001111000000;
		15'h2109: char_row_bitmap <= 16'b0000001111000000;
		15'h210a: char_row_bitmap <= 16'b0000001111000000;
		15'h210b: char_row_bitmap <= 16'b0000001111000000;
		15'h210c: char_row_bitmap <= 16'b0000001111000000;
		15'h210d: char_row_bitmap <= 16'b0000001111000000;
		15'h210e: char_row_bitmap <= 16'b0000001111000000;
		15'h210f: char_row_bitmap <= 16'b0000001111000000;
		15'h2110: char_row_bitmap <= 16'b0000001111000000;
		15'h2111: char_row_bitmap <= 16'b0000001111000000;
		15'h2112: char_row_bitmap <= 16'b0000001111000000;
		15'h2113: char_row_bitmap <= 16'b0000001111000000;
		15'h2114: char_row_bitmap <= 16'b0000001111111111;
		15'h2115: char_row_bitmap <= 16'b0000001111111111;
		15'h2116: char_row_bitmap <= 16'b0000001111111111;
		15'h2117: char_row_bitmap <= 16'b0000001111111111;
		15'h2118: char_row_bitmap <= 16'b0000001111000000;
		15'h2119: char_row_bitmap <= 16'b0000001111000000;
		15'h211a: char_row_bitmap <= 16'b0000001111000000;
		15'h211b: char_row_bitmap <= 16'b0000001111000000;
		15'h211c: char_row_bitmap <= 16'b0000001111000000;
		15'h211d: char_row_bitmap <= 16'b0000001111000000;
		15'h211e: char_row_bitmap <= 16'b0000001111000000;
		15'h211f: char_row_bitmap <= 16'b0000001111000000;
		15'h2120: char_row_bitmap <= 16'b0000000000000000;
		15'h2121: char_row_bitmap <= 16'b0000000000000000;
		15'h2122: char_row_bitmap <= 16'b0000000000000000;
		15'h2123: char_row_bitmap <= 16'b0000000000000000;
		15'h2124: char_row_bitmap <= 16'b0000000000000000;
		15'h2125: char_row_bitmap <= 16'b0000000000000000;
		15'h2126: char_row_bitmap <= 16'b0000000000000000;
		15'h2127: char_row_bitmap <= 16'b0000000000000000;
		15'h2128: char_row_bitmap <= 16'b1111111111000000;
		15'h2129: char_row_bitmap <= 16'b1111111111000000;
		15'h212a: char_row_bitmap <= 16'b1111111111000000;
		15'h212b: char_row_bitmap <= 16'b1111111111000000;
		15'h212c: char_row_bitmap <= 16'b0000000000000000;
		15'h212d: char_row_bitmap <= 16'b0000000000000000;
		15'h212e: char_row_bitmap <= 16'b0000000000000000;
		15'h212f: char_row_bitmap <= 16'b0000000000000000;
		15'h2130: char_row_bitmap <= 16'b0000000000000000;
		15'h2131: char_row_bitmap <= 16'b0000000000000000;
		15'h2132: char_row_bitmap <= 16'b0000000000000000;
		15'h2133: char_row_bitmap <= 16'b0000000000000000;
		15'h2134: char_row_bitmap <= 16'b0000001111000000;
		15'h2135: char_row_bitmap <= 16'b0000001111000000;
		15'h2136: char_row_bitmap <= 16'b0000001111000000;
		15'h2137: char_row_bitmap <= 16'b0000001111000000;
		15'h2138: char_row_bitmap <= 16'b0000001111000000;
		15'h2139: char_row_bitmap <= 16'b0000001111000000;
		15'h213a: char_row_bitmap <= 16'b0000001111000000;
		15'h213b: char_row_bitmap <= 16'b0000001111000000;
		15'h213c: char_row_bitmap <= 16'b1111111111000000;
		15'h213d: char_row_bitmap <= 16'b1111111111000000;
		15'h213e: char_row_bitmap <= 16'b1111111111000000;
		15'h213f: char_row_bitmap <= 16'b1111111111000000;
		15'h2140: char_row_bitmap <= 16'b0000000000000000;
		15'h2141: char_row_bitmap <= 16'b0000000000000000;
		15'h2142: char_row_bitmap <= 16'b0000000000000000;
		15'h2143: char_row_bitmap <= 16'b0000000000000000;
		15'h2144: char_row_bitmap <= 16'b0000000000000000;
		15'h2145: char_row_bitmap <= 16'b0000000000000000;
		15'h2146: char_row_bitmap <= 16'b0000000000000000;
		15'h2147: char_row_bitmap <= 16'b0000000000000000;
		15'h2148: char_row_bitmap <= 16'b0000000000000000;
		15'h2149: char_row_bitmap <= 16'b0000000000000000;
		15'h214a: char_row_bitmap <= 16'b0000000000000000;
		15'h214b: char_row_bitmap <= 16'b0000000000000000;
		15'h214c: char_row_bitmap <= 16'b0000000000000000;
		15'h214d: char_row_bitmap <= 16'b0000000000000000;
		15'h214e: char_row_bitmap <= 16'b0000000000000000;
		15'h214f: char_row_bitmap <= 16'b0000000000000000;
		15'h2150: char_row_bitmap <= 16'b1111111111111111;
		15'h2151: char_row_bitmap <= 16'b1111111111111111;
		15'h2152: char_row_bitmap <= 16'b1111111111111111;
		15'h2153: char_row_bitmap <= 16'b1111111111111111;
		15'h2154: char_row_bitmap <= 16'b0000000000000000;
		15'h2155: char_row_bitmap <= 16'b0000000000000000;
		15'h2156: char_row_bitmap <= 16'b0000000000000000;
		15'h2157: char_row_bitmap <= 16'b0000000000000000;
		15'h2158: char_row_bitmap <= 16'b0000000000000000;
		15'h2159: char_row_bitmap <= 16'b0000000000000000;
		15'h215a: char_row_bitmap <= 16'b0000000000000000;
		15'h215b: char_row_bitmap <= 16'b0000000000000000;
		15'h215c: char_row_bitmap <= 16'b0000001111000000;
		15'h215d: char_row_bitmap <= 16'b0000001111000000;
		15'h215e: char_row_bitmap <= 16'b0000001111000000;
		15'h215f: char_row_bitmap <= 16'b0000001111000000;
		15'h2160: char_row_bitmap <= 16'b0000001111000000;
		15'h2161: char_row_bitmap <= 16'b0000001111000000;
		15'h2162: char_row_bitmap <= 16'b0000001111000000;
		15'h2163: char_row_bitmap <= 16'b0000001111000000;
		15'h2164: char_row_bitmap <= 16'b1111111111111111;
		15'h2165: char_row_bitmap <= 16'b1111111111111111;
		15'h2166: char_row_bitmap <= 16'b1111111111111111;
		15'h2167: char_row_bitmap <= 16'b1111111111111111;
		15'h2168: char_row_bitmap <= 16'b0000000000000000;
		15'h2169: char_row_bitmap <= 16'b0000000000000000;
		15'h216a: char_row_bitmap <= 16'b0000000000000000;
		15'h216b: char_row_bitmap <= 16'b0000000000000000;
		15'h216c: char_row_bitmap <= 16'b0000000000000000;
		15'h216d: char_row_bitmap <= 16'b0000000000000000;
		15'h216e: char_row_bitmap <= 16'b0000000000000000;
		15'h216f: char_row_bitmap <= 16'b0000000000000000;
		15'h2170: char_row_bitmap <= 16'b0000000000000000;
		15'h2171: char_row_bitmap <= 16'b0000000000000000;
		15'h2172: char_row_bitmap <= 16'b0000000000000000;
		15'h2173: char_row_bitmap <= 16'b0000000000000000;
		15'h2174: char_row_bitmap <= 16'b0000000000000000;
		15'h2175: char_row_bitmap <= 16'b0000000000000000;
		15'h2176: char_row_bitmap <= 16'b0000000000000000;
		15'h2177: char_row_bitmap <= 16'b0000000000000000;
		15'h2178: char_row_bitmap <= 16'b1111111111000000;
		15'h2179: char_row_bitmap <= 16'b1111111111000000;
		15'h217a: char_row_bitmap <= 16'b1111111111000000;
		15'h217b: char_row_bitmap <= 16'b1111111111000000;
		15'h217c: char_row_bitmap <= 16'b0000001111000000;
		15'h217d: char_row_bitmap <= 16'b0000001111000000;
		15'h217e: char_row_bitmap <= 16'b0000001111000000;
		15'h217f: char_row_bitmap <= 16'b0000001111000000;
		15'h2180: char_row_bitmap <= 16'b0000001111000000;
		15'h2181: char_row_bitmap <= 16'b0000001111000000;
		15'h2182: char_row_bitmap <= 16'b0000001111000000;
		15'h2183: char_row_bitmap <= 16'b0000001111000000;
		15'h2184: char_row_bitmap <= 16'b0000001111000000;
		15'h2185: char_row_bitmap <= 16'b0000001111000000;
		15'h2186: char_row_bitmap <= 16'b0000001111000000;
		15'h2187: char_row_bitmap <= 16'b0000001111000000;
		15'h2188: char_row_bitmap <= 16'b0000001111000000;
		15'h2189: char_row_bitmap <= 16'b0000001111000000;
		15'h218a: char_row_bitmap <= 16'b0000001111000000;
		15'h218b: char_row_bitmap <= 16'b0000001111000000;
		15'h218c: char_row_bitmap <= 16'b1111111111000000;
		15'h218d: char_row_bitmap <= 16'b1111111111000000;
		15'h218e: char_row_bitmap <= 16'b1111111111000000;
		15'h218f: char_row_bitmap <= 16'b1111111111000000;
		15'h2190: char_row_bitmap <= 16'b0000001111000000;
		15'h2191: char_row_bitmap <= 16'b0000001111000000;
		15'h2192: char_row_bitmap <= 16'b0000001111000000;
		15'h2193: char_row_bitmap <= 16'b0000001111000000;
		15'h2194: char_row_bitmap <= 16'b0000001111000000;
		15'h2195: char_row_bitmap <= 16'b0000001111000000;
		15'h2196: char_row_bitmap <= 16'b0000001111000000;
		15'h2197: char_row_bitmap <= 16'b0000001111000000;
		15'h2198: char_row_bitmap <= 16'b0000000000000000;
		15'h2199: char_row_bitmap <= 16'b0000000000000000;
		15'h219a: char_row_bitmap <= 16'b0000000000000000;
		15'h219b: char_row_bitmap <= 16'b0000000000000000;
		15'h219c: char_row_bitmap <= 16'b0000000000000000;
		15'h219d: char_row_bitmap <= 16'b0000000000000000;
		15'h219e: char_row_bitmap <= 16'b0000000000000000;
		15'h219f: char_row_bitmap <= 16'b0000000000000000;
		15'h21a0: char_row_bitmap <= 16'b1111111111111111;
		15'h21a1: char_row_bitmap <= 16'b1111111111111111;
		15'h21a2: char_row_bitmap <= 16'b1111111111111111;
		15'h21a3: char_row_bitmap <= 16'b1111111111111111;
		15'h21a4: char_row_bitmap <= 16'b0000001111000000;
		15'h21a5: char_row_bitmap <= 16'b0000001111000000;
		15'h21a6: char_row_bitmap <= 16'b0000001111000000;
		15'h21a7: char_row_bitmap <= 16'b0000001111000000;
		15'h21a8: char_row_bitmap <= 16'b0000001111000000;
		15'h21a9: char_row_bitmap <= 16'b0000001111000000;
		15'h21aa: char_row_bitmap <= 16'b0000001111000000;
		15'h21ab: char_row_bitmap <= 16'b0000001111000000;
		15'h21ac: char_row_bitmap <= 16'b0000001111000000;
		15'h21ad: char_row_bitmap <= 16'b0000001111000000;
		15'h21ae: char_row_bitmap <= 16'b0000001111000000;
		15'h21af: char_row_bitmap <= 16'b0000001111000000;
		15'h21b0: char_row_bitmap <= 16'b0000001111000000;
		15'h21b1: char_row_bitmap <= 16'b0000001111000000;
		15'h21b2: char_row_bitmap <= 16'b0000001111000000;
		15'h21b3: char_row_bitmap <= 16'b0000001111000000;
		15'h21b4: char_row_bitmap <= 16'b1111111111111111;
		15'h21b5: char_row_bitmap <= 16'b1111111111111111;
		15'h21b6: char_row_bitmap <= 16'b1111111111111111;
		15'h21b7: char_row_bitmap <= 16'b1111111111111111;
		15'h21b8: char_row_bitmap <= 16'b0000001111000000;
		15'h21b9: char_row_bitmap <= 16'b0000001111000000;
		15'h21ba: char_row_bitmap <= 16'b0000001111000000;
		15'h21bb: char_row_bitmap <= 16'b0000001111000000;
		15'h21bc: char_row_bitmap <= 16'b0000001111000000;
		15'h21bd: char_row_bitmap <= 16'b0000001111000000;
		15'h21be: char_row_bitmap <= 16'b0000001111000000;
		15'h21bf: char_row_bitmap <= 16'b0000001111000000;
		15'h21c0: char_row_bitmap <= 16'b0000001001000000;
		15'h21c1: char_row_bitmap <= 16'b0000001001000000;
		15'h21c2: char_row_bitmap <= 16'b0000001001000000;
		15'h21c3: char_row_bitmap <= 16'b0000000000000000;
		15'h21c4: char_row_bitmap <= 16'b0000000000000000;
		15'h21c5: char_row_bitmap <= 16'b0000001001000000;
		15'h21c6: char_row_bitmap <= 16'b0000001001000000;
		15'h21c7: char_row_bitmap <= 16'b0000001001000000;
		15'h21c8: char_row_bitmap <= 16'b0000001001000000;
		15'h21c9: char_row_bitmap <= 16'b0000000000000000;
		15'h21ca: char_row_bitmap <= 16'b0000000000000000;
		15'h21cb: char_row_bitmap <= 16'b0000001001000000;
		15'h21cc: char_row_bitmap <= 16'b0000001001000000;
		15'h21cd: char_row_bitmap <= 16'b0000001001000000;
		15'h21ce: char_row_bitmap <= 16'b0000001001000000;
		15'h21cf: char_row_bitmap <= 16'b0000000000000000;
		15'h21d0: char_row_bitmap <= 16'b0000000000000000;
		15'h21d1: char_row_bitmap <= 16'b0000001001000000;
		15'h21d2: char_row_bitmap <= 16'b0000001001000000;
		15'h21d3: char_row_bitmap <= 16'b0000001001000000;
		15'h21d4: char_row_bitmap <= 16'b0000000110000000;
		15'h21d5: char_row_bitmap <= 16'b0000000110000000;
		15'h21d6: char_row_bitmap <= 16'b0000000110000000;
		15'h21d7: char_row_bitmap <= 16'b0000000000000000;
		15'h21d8: char_row_bitmap <= 16'b0000000000000000;
		15'h21d9: char_row_bitmap <= 16'b0000000110000000;
		15'h21da: char_row_bitmap <= 16'b0000000110000000;
		15'h21db: char_row_bitmap <= 16'b0000000110000000;
		15'h21dc: char_row_bitmap <= 16'b0000000110000000;
		15'h21dd: char_row_bitmap <= 16'b0000000000000000;
		15'h21de: char_row_bitmap <= 16'b0000000000000000;
		15'h21df: char_row_bitmap <= 16'b0000000110000000;
		15'h21e0: char_row_bitmap <= 16'b0000000110000000;
		15'h21e1: char_row_bitmap <= 16'b0000000110000000;
		15'h21e2: char_row_bitmap <= 16'b0000000110000000;
		15'h21e3: char_row_bitmap <= 16'b0000000000000000;
		15'h21e4: char_row_bitmap <= 16'b0000000000000000;
		15'h21e5: char_row_bitmap <= 16'b0000000110000000;
		15'h21e6: char_row_bitmap <= 16'b0000000110000000;
		15'h21e7: char_row_bitmap <= 16'b0000000110000000;
		15'h21e8: char_row_bitmap <= 16'b0000001111000000;
		15'h21e9: char_row_bitmap <= 16'b0000001111000000;
		15'h21ea: char_row_bitmap <= 16'b0000001111000000;
		15'h21eb: char_row_bitmap <= 16'b0000000000000000;
		15'h21ec: char_row_bitmap <= 16'b0000000000000000;
		15'h21ed: char_row_bitmap <= 16'b0000001111000000;
		15'h21ee: char_row_bitmap <= 16'b0000001111000000;
		15'h21ef: char_row_bitmap <= 16'b0000001111000000;
		15'h21f0: char_row_bitmap <= 16'b0000001111000000;
		15'h21f1: char_row_bitmap <= 16'b0000000000000000;
		15'h21f2: char_row_bitmap <= 16'b0000000000000000;
		15'h21f3: char_row_bitmap <= 16'b0000001111000000;
		15'h21f4: char_row_bitmap <= 16'b0000001111000000;
		15'h21f5: char_row_bitmap <= 16'b0000001111000000;
		15'h21f6: char_row_bitmap <= 16'b0000001111000000;
		15'h21f7: char_row_bitmap <= 16'b0000000000000000;
		15'h21f8: char_row_bitmap <= 16'b0000000000000000;
		15'h21f9: char_row_bitmap <= 16'b0000001111000000;
		15'h21fa: char_row_bitmap <= 16'b0000001111000000;
		15'h21fb: char_row_bitmap <= 16'b0000001111000000;
		15'h21fc: char_row_bitmap <= 16'b0000000000000000;
		15'h21fd: char_row_bitmap <= 16'b0000000000000000;
		15'h21fe: char_row_bitmap <= 16'b0000000000000000;
		15'h21ff: char_row_bitmap <= 16'b0000000000000000;
		15'h2200: char_row_bitmap <= 16'b0000000000000000;
		15'h2201: char_row_bitmap <= 16'b0000000000000000;
		15'h2202: char_row_bitmap <= 16'b0000000000000000;
		15'h2203: char_row_bitmap <= 16'b0000000000000000;
		15'h2204: char_row_bitmap <= 16'b1100111001110011;
		15'h2205: char_row_bitmap <= 16'b0000000000000000;
		15'h2206: char_row_bitmap <= 16'b0000000000000000;
		15'h2207: char_row_bitmap <= 16'b1100111001110011;
		15'h2208: char_row_bitmap <= 16'b0000000000000000;
		15'h2209: char_row_bitmap <= 16'b0000000000000000;
		15'h220a: char_row_bitmap <= 16'b0000000000000000;
		15'h220b: char_row_bitmap <= 16'b0000000000000000;
		15'h220c: char_row_bitmap <= 16'b0000000000000000;
		15'h220d: char_row_bitmap <= 16'b0000000000000000;
		15'h220e: char_row_bitmap <= 16'b0000000000000000;
		15'h220f: char_row_bitmap <= 16'b0000000000000000;
		15'h2210: char_row_bitmap <= 16'b0000000000000000;
		15'h2211: char_row_bitmap <= 16'b0000000000000000;
		15'h2212: char_row_bitmap <= 16'b0000000000000000;
		15'h2213: char_row_bitmap <= 16'b0000000000000000;
		15'h2214: char_row_bitmap <= 16'b0000000000000000;
		15'h2215: char_row_bitmap <= 16'b0000000000000000;
		15'h2216: char_row_bitmap <= 16'b0000000000000000;
		15'h2217: char_row_bitmap <= 16'b0000000000000000;
		15'h2218: char_row_bitmap <= 16'b0000000000000000;
		15'h2219: char_row_bitmap <= 16'b1100111001110011;
		15'h221a: char_row_bitmap <= 16'b1100111001110011;
		15'h221b: char_row_bitmap <= 16'b0000000000000000;
		15'h221c: char_row_bitmap <= 16'b0000000000000000;
		15'h221d: char_row_bitmap <= 16'b0000000000000000;
		15'h221e: char_row_bitmap <= 16'b0000000000000000;
		15'h221f: char_row_bitmap <= 16'b0000000000000000;
		15'h2220: char_row_bitmap <= 16'b0000000000000000;
		15'h2221: char_row_bitmap <= 16'b0000000000000000;
		15'h2222: char_row_bitmap <= 16'b0000000000000000;
		15'h2223: char_row_bitmap <= 16'b0000000000000000;
		15'h2224: char_row_bitmap <= 16'b0000000000000000;
		15'h2225: char_row_bitmap <= 16'b0000000000000000;
		15'h2226: char_row_bitmap <= 16'b0000000000000000;
		15'h2227: char_row_bitmap <= 16'b0000000000000000;
		15'h2228: char_row_bitmap <= 16'b0000000000000000;
		15'h2229: char_row_bitmap <= 16'b0000000000000000;
		15'h222a: char_row_bitmap <= 16'b0000000000000000;
		15'h222b: char_row_bitmap <= 16'b0000000000000000;
		15'h222c: char_row_bitmap <= 16'b1100111001110011;
		15'h222d: char_row_bitmap <= 16'b1100111001110011;
		15'h222e: char_row_bitmap <= 16'b1100111001110011;
		15'h222f: char_row_bitmap <= 16'b1100111001110011;
		15'h2230: char_row_bitmap <= 16'b0000000000000000;
		15'h2231: char_row_bitmap <= 16'b0000000000000000;
		15'h2232: char_row_bitmap <= 16'b0000000000000000;
		15'h2233: char_row_bitmap <= 16'b0000000000000000;
		15'h2234: char_row_bitmap <= 16'b0000000000000000;
		15'h2235: char_row_bitmap <= 16'b0000000000000000;
		15'h2236: char_row_bitmap <= 16'b0000000000000000;
		15'h2237: char_row_bitmap <= 16'b0000000000000000;
		15'h2238: char_row_bitmap <= 16'b0000001001000000;
		15'h2239: char_row_bitmap <= 16'b0000001001000000;
		15'h223a: char_row_bitmap <= 16'b0000001001000000;
		15'h223b: char_row_bitmap <= 16'b0000001001000000;
		15'h223c: char_row_bitmap <= 16'b0000001001000000;
		15'h223d: char_row_bitmap <= 16'b0000001001000000;
		15'h223e: char_row_bitmap <= 16'b0000001001000000;
		15'h223f: char_row_bitmap <= 16'b0000001001000000;
		15'h2240: char_row_bitmap <= 16'b0000001001000000;
		15'h2241: char_row_bitmap <= 16'b0000001001111111;
		15'h2242: char_row_bitmap <= 16'b0000001001111111;
		15'h2243: char_row_bitmap <= 16'b0000001001000000;
		15'h2244: char_row_bitmap <= 16'b0000001001000000;
		15'h2245: char_row_bitmap <= 16'b0000001001000000;
		15'h2246: char_row_bitmap <= 16'b0000001001000000;
		15'h2247: char_row_bitmap <= 16'b0000001001000000;
		15'h2248: char_row_bitmap <= 16'b0000001001000000;
		15'h2249: char_row_bitmap <= 16'b0000001001000000;
		15'h224a: char_row_bitmap <= 16'b0000001001000000;
		15'h224b: char_row_bitmap <= 16'b0000001001000000;
		15'h224c: char_row_bitmap <= 16'b0000001001000000;
		15'h224d: char_row_bitmap <= 16'b0000001001000000;
		15'h224e: char_row_bitmap <= 16'b0000001001000000;
		15'h224f: char_row_bitmap <= 16'b0000001001000000;
		15'h2250: char_row_bitmap <= 16'b0000001001000000;
		15'h2251: char_row_bitmap <= 16'b0000001001000000;
		15'h2252: char_row_bitmap <= 16'b0000001001000000;
		15'h2253: char_row_bitmap <= 16'b0000001001000000;
		15'h2254: char_row_bitmap <= 16'b0000001001000000;
		15'h2255: char_row_bitmap <= 16'b1111111001000000;
		15'h2256: char_row_bitmap <= 16'b1111111001000000;
		15'h2257: char_row_bitmap <= 16'b0000001001000000;
		15'h2258: char_row_bitmap <= 16'b0000001001000000;
		15'h2259: char_row_bitmap <= 16'b0000001001000000;
		15'h225a: char_row_bitmap <= 16'b0000001001000000;
		15'h225b: char_row_bitmap <= 16'b0000001001000000;
		15'h225c: char_row_bitmap <= 16'b0000001001000000;
		15'h225d: char_row_bitmap <= 16'b0000001001000000;
		15'h225e: char_row_bitmap <= 16'b0000001001000000;
		15'h225f: char_row_bitmap <= 16'b0000001001000000;
		15'h2260: char_row_bitmap <= 16'b0000000110000000;
		15'h2261: char_row_bitmap <= 16'b0000000110000000;
		15'h2262: char_row_bitmap <= 16'b0000000110000000;
		15'h2263: char_row_bitmap <= 16'b0000000110000000;
		15'h2264: char_row_bitmap <= 16'b0000000110000000;
		15'h2265: char_row_bitmap <= 16'b0000000110000000;
		15'h2266: char_row_bitmap <= 16'b0000000110000000;
		15'h2267: char_row_bitmap <= 16'b0000000110000000;
		15'h2268: char_row_bitmap <= 16'b1111111111111111;
		15'h2269: char_row_bitmap <= 16'b0000000000000000;
		15'h226a: char_row_bitmap <= 16'b0000000000000000;
		15'h226b: char_row_bitmap <= 16'b1111111111111111;
		15'h226c: char_row_bitmap <= 16'b0000000000000000;
		15'h226d: char_row_bitmap <= 16'b0000000000000000;
		15'h226e: char_row_bitmap <= 16'b0000000000000000;
		15'h226f: char_row_bitmap <= 16'b0000000000000000;
		15'h2270: char_row_bitmap <= 16'b0000000000000000;
		15'h2271: char_row_bitmap <= 16'b0000000000000000;
		15'h2272: char_row_bitmap <= 16'b0000000000000000;
		15'h2273: char_row_bitmap <= 16'b0000000000000000;
		15'h2274: char_row_bitmap <= 16'b0000000000000000;
		15'h2275: char_row_bitmap <= 16'b0000000000000000;
		15'h2276: char_row_bitmap <= 16'b0000000000000000;
		15'h2277: char_row_bitmap <= 16'b0000000000000000;
		15'h2278: char_row_bitmap <= 16'b0000000000000000;
		15'h2279: char_row_bitmap <= 16'b0000000000000000;
		15'h227a: char_row_bitmap <= 16'b0000000000000000;
		15'h227b: char_row_bitmap <= 16'b0000000000000000;
		15'h227c: char_row_bitmap <= 16'b1111111111111111;
		15'h227d: char_row_bitmap <= 16'b0000000000000000;
		15'h227e: char_row_bitmap <= 16'b0000000000000000;
		15'h227f: char_row_bitmap <= 16'b1111111111111111;
		15'h2280: char_row_bitmap <= 16'b0000000110000000;
		15'h2281: char_row_bitmap <= 16'b0000000110000000;
		15'h2282: char_row_bitmap <= 16'b0000000110000000;
		15'h2283: char_row_bitmap <= 16'b0000000110000000;
		15'h2284: char_row_bitmap <= 16'b0000000110000000;
		15'h2285: char_row_bitmap <= 16'b0000000110000000;
		15'h2286: char_row_bitmap <= 16'b0000000110000000;
		15'h2287: char_row_bitmap <= 16'b0000000110000000;
		15'h2288: char_row_bitmap <= 16'b0000000110000000;
		15'h2289: char_row_bitmap <= 16'b0000000110000000;
		15'h228a: char_row_bitmap <= 16'b0000000110000000;
		15'h228b: char_row_bitmap <= 16'b0000000110000000;
		15'h228c: char_row_bitmap <= 16'b0000000110000000;
		15'h228d: char_row_bitmap <= 16'b0000000110000000;
		15'h228e: char_row_bitmap <= 16'b0000000110000000;
		15'h228f: char_row_bitmap <= 16'b0000000110000000;
		15'h2290: char_row_bitmap <= 16'b1111111111111111;
		15'h2291: char_row_bitmap <= 16'b1111111111111111;
		15'h2292: char_row_bitmap <= 16'b1111111111111111;
		15'h2293: char_row_bitmap <= 16'b1111111111111111;
		15'h2294: char_row_bitmap <= 16'b0000001111000000;
		15'h2295: char_row_bitmap <= 16'b0000001111000000;
		15'h2296: char_row_bitmap <= 16'b0000001111000000;
		15'h2297: char_row_bitmap <= 16'b0000001111000000;
		15'h2298: char_row_bitmap <= 16'b0000001111000000;
		15'h2299: char_row_bitmap <= 16'b0000001111000000;
		15'h229a: char_row_bitmap <= 16'b0000001111000000;
		15'h229b: char_row_bitmap <= 16'b0000001111000000;
		15'h229c: char_row_bitmap <= 16'b0000001111000000;
		15'h229d: char_row_bitmap <= 16'b0000001111000000;
		15'h229e: char_row_bitmap <= 16'b0000001111000000;
		15'h229f: char_row_bitmap <= 16'b0000001111000000;
		15'h22a0: char_row_bitmap <= 16'b0000001111000000;
		15'h22a1: char_row_bitmap <= 16'b0000001111000000;
		15'h22a2: char_row_bitmap <= 16'b0000001111000000;
		15'h22a3: char_row_bitmap <= 16'b0000001111000000;
		15'h22a4: char_row_bitmap <= 16'b0000001111111111;
		15'h22a5: char_row_bitmap <= 16'b1111111111111111;
		15'h22a6: char_row_bitmap <= 16'b1111111111111111;
		15'h22a7: char_row_bitmap <= 16'b0000001111111111;
		15'h22a8: char_row_bitmap <= 16'b0000001111000000;
		15'h22a9: char_row_bitmap <= 16'b0000001111000000;
		15'h22aa: char_row_bitmap <= 16'b0000001111000000;
		15'h22ab: char_row_bitmap <= 16'b0000001111000000;
		15'h22ac: char_row_bitmap <= 16'b0000001111000000;
		15'h22ad: char_row_bitmap <= 16'b0000001111000000;
		15'h22ae: char_row_bitmap <= 16'b0000001111000000;
		15'h22af: char_row_bitmap <= 16'b0000001111000000;
		15'h22b0: char_row_bitmap <= 16'b0000001111000000;
		15'h22b1: char_row_bitmap <= 16'b0000001111000000;
		15'h22b2: char_row_bitmap <= 16'b0000001111000000;
		15'h22b3: char_row_bitmap <= 16'b0000001111000000;
		15'h22b4: char_row_bitmap <= 16'b0000001111000000;
		15'h22b5: char_row_bitmap <= 16'b0000001111000000;
		15'h22b6: char_row_bitmap <= 16'b0000001111000000;
		15'h22b7: char_row_bitmap <= 16'b0000001111000000;
		15'h22b8: char_row_bitmap <= 16'b1111111111111111;
		15'h22b9: char_row_bitmap <= 16'b1111111111111111;
		15'h22ba: char_row_bitmap <= 16'b1111111111111111;
		15'h22bb: char_row_bitmap <= 16'b1111111111111111;
		15'h22bc: char_row_bitmap <= 16'b0000000110000000;
		15'h22bd: char_row_bitmap <= 16'b0000000110000000;
		15'h22be: char_row_bitmap <= 16'b0000000110000000;
		15'h22bf: char_row_bitmap <= 16'b0000000110000000;
		15'h22c0: char_row_bitmap <= 16'b0000000110000000;
		15'h22c1: char_row_bitmap <= 16'b0000000110000000;
		15'h22c2: char_row_bitmap <= 16'b0000000110000000;
		15'h22c3: char_row_bitmap <= 16'b0000000110000000;
		15'h22c4: char_row_bitmap <= 16'b0000001111000000;
		15'h22c5: char_row_bitmap <= 16'b0000001111000000;
		15'h22c6: char_row_bitmap <= 16'b0000001111000000;
		15'h22c7: char_row_bitmap <= 16'b0000001111000000;
		15'h22c8: char_row_bitmap <= 16'b0000001111000000;
		15'h22c9: char_row_bitmap <= 16'b0000001111000000;
		15'h22ca: char_row_bitmap <= 16'b0000001111000000;
		15'h22cb: char_row_bitmap <= 16'b0000001111000000;
		15'h22cc: char_row_bitmap <= 16'b1111111111000000;
		15'h22cd: char_row_bitmap <= 16'b1111111111111111;
		15'h22ce: char_row_bitmap <= 16'b1111111111111111;
		15'h22cf: char_row_bitmap <= 16'b1111111111000000;
		15'h22d0: char_row_bitmap <= 16'b0000001111000000;
		15'h22d1: char_row_bitmap <= 16'b0000001111000000;
		15'h22d2: char_row_bitmap <= 16'b0000001111000000;
		15'h22d3: char_row_bitmap <= 16'b0000001111000000;
		15'h22d4: char_row_bitmap <= 16'b0000001111000000;
		15'h22d5: char_row_bitmap <= 16'b0000001111000000;
		15'h22d6: char_row_bitmap <= 16'b0000001111000000;
		15'h22d7: char_row_bitmap <= 16'b0000001111000000;
		15'h22d8: char_row_bitmap <= 16'b0000000110000000;
		15'h22d9: char_row_bitmap <= 16'b0000000110000000;
		15'h22da: char_row_bitmap <= 16'b0000000110000000;
		15'h22db: char_row_bitmap <= 16'b0000000110000000;
		15'h22dc: char_row_bitmap <= 16'b0000000110000000;
		15'h22dd: char_row_bitmap <= 16'b0000000110000000;
		15'h22de: char_row_bitmap <= 16'b0000000110000000;
		15'h22df: char_row_bitmap <= 16'b0000000110000000;
		15'h22e0: char_row_bitmap <= 16'b1111111111111111;
		15'h22e1: char_row_bitmap <= 16'b1111111111111111;
		15'h22e2: char_row_bitmap <= 16'b1111111111111111;
		15'h22e3: char_row_bitmap <= 16'b1111111111111111;
		15'h22e4: char_row_bitmap <= 16'b0000000110000000;
		15'h22e5: char_row_bitmap <= 16'b0000000110000000;
		15'h22e6: char_row_bitmap <= 16'b0000000110000000;
		15'h22e7: char_row_bitmap <= 16'b0000000110000000;
		15'h22e8: char_row_bitmap <= 16'b0000000110000000;
		15'h22e9: char_row_bitmap <= 16'b0000000110000000;
		15'h22ea: char_row_bitmap <= 16'b0000000110000000;
		15'h22eb: char_row_bitmap <= 16'b0000000110000000;
		15'h22ec: char_row_bitmap <= 16'b0000001111000000;
		15'h22ed: char_row_bitmap <= 16'b0000001111000000;
		15'h22ee: char_row_bitmap <= 16'b0000001111000000;
		15'h22ef: char_row_bitmap <= 16'b0000001111000000;
		15'h22f0: char_row_bitmap <= 16'b0000001111000000;
		15'h22f1: char_row_bitmap <= 16'b0000001111000000;
		15'h22f2: char_row_bitmap <= 16'b0000001111000000;
		15'h22f3: char_row_bitmap <= 16'b0000001111000000;
		15'h22f4: char_row_bitmap <= 16'b0000001111000000;
		15'h22f5: char_row_bitmap <= 16'b1111111111111111;
		15'h22f6: char_row_bitmap <= 16'b1111111111111111;
		15'h22f7: char_row_bitmap <= 16'b0000001111000000;
		15'h22f8: char_row_bitmap <= 16'b0000001111000000;
		15'h22f9: char_row_bitmap <= 16'b0000001111000000;
		15'h22fa: char_row_bitmap <= 16'b0000001111000000;
		15'h22fb: char_row_bitmap <= 16'b0000001111000000;
		15'h22fc: char_row_bitmap <= 16'b0000001111000000;
		15'h22fd: char_row_bitmap <= 16'b0000001111000000;
		15'h22fe: char_row_bitmap <= 16'b0000001111000000;
		15'h22ff: char_row_bitmap <= 16'b0000001111000000;
		15'h2300: char_row_bitmap <= 16'b0000001111000000;
		15'h2301: char_row_bitmap <= 16'b0000001111000000;
		15'h2302: char_row_bitmap <= 16'b0000001111000000;
		15'h2303: char_row_bitmap <= 16'b0000001111000000;
		15'h2304: char_row_bitmap <= 16'b0000001111000000;
		15'h2305: char_row_bitmap <= 16'b0000001111000000;
		15'h2306: char_row_bitmap <= 16'b0000001111000000;
		15'h2307: char_row_bitmap <= 16'b0000001111000000;
		15'h2308: char_row_bitmap <= 16'b0000001111000000;
		15'h2309: char_row_bitmap <= 16'b0000001111111111;
		15'h230a: char_row_bitmap <= 16'b0000001111111111;
		15'h230b: char_row_bitmap <= 16'b0000000000000000;
		15'h230c: char_row_bitmap <= 16'b0000000000000000;
		15'h230d: char_row_bitmap <= 16'b0000000000000000;
		15'h230e: char_row_bitmap <= 16'b0000000000000000;
		15'h230f: char_row_bitmap <= 16'b0000000000000000;
		15'h2310: char_row_bitmap <= 16'b0000000000000000;
		15'h2311: char_row_bitmap <= 16'b0000000000000000;
		15'h2312: char_row_bitmap <= 16'b0000000000000000;
		15'h2313: char_row_bitmap <= 16'b0000000000000000;
		15'h2314: char_row_bitmap <= 16'b0000000110000000;
		15'h2315: char_row_bitmap <= 16'b0000000110000000;
		15'h2316: char_row_bitmap <= 16'b0000000110000000;
		15'h2317: char_row_bitmap <= 16'b0000000110000000;
		15'h2318: char_row_bitmap <= 16'b0000000110000000;
		15'h2319: char_row_bitmap <= 16'b0000000110000000;
		15'h231a: char_row_bitmap <= 16'b0000000110000000;
		15'h231b: char_row_bitmap <= 16'b0000000110000000;
		15'h231c: char_row_bitmap <= 16'b0000000111111111;
		15'h231d: char_row_bitmap <= 16'b0000000111111111;
		15'h231e: char_row_bitmap <= 16'b0000000111111111;
		15'h231f: char_row_bitmap <= 16'b0000000111111111;
		15'h2320: char_row_bitmap <= 16'b0000000000000000;
		15'h2321: char_row_bitmap <= 16'b0000000000000000;
		15'h2322: char_row_bitmap <= 16'b0000000000000000;
		15'h2323: char_row_bitmap <= 16'b0000000000000000;
		15'h2324: char_row_bitmap <= 16'b0000000000000000;
		15'h2325: char_row_bitmap <= 16'b0000000000000000;
		15'h2326: char_row_bitmap <= 16'b0000000000000000;
		15'h2327: char_row_bitmap <= 16'b0000000000000000;
		15'h2328: char_row_bitmap <= 16'b0000000000000000;
		15'h2329: char_row_bitmap <= 16'b0000000000000000;
		15'h232a: char_row_bitmap <= 16'b0000000000000000;
		15'h232b: char_row_bitmap <= 16'b0000000000000000;
		15'h232c: char_row_bitmap <= 16'b0000000000000000;
		15'h232d: char_row_bitmap <= 16'b0000000000000000;
		15'h232e: char_row_bitmap <= 16'b0000000000000000;
		15'h232f: char_row_bitmap <= 16'b0000000000000000;
		15'h2330: char_row_bitmap <= 16'b0000000000000000;
		15'h2331: char_row_bitmap <= 16'b0000001111111111;
		15'h2332: char_row_bitmap <= 16'b0000001111111111;
		15'h2333: char_row_bitmap <= 16'b0000001111000000;
		15'h2334: char_row_bitmap <= 16'b0000001111000000;
		15'h2335: char_row_bitmap <= 16'b0000001111000000;
		15'h2336: char_row_bitmap <= 16'b0000001111000000;
		15'h2337: char_row_bitmap <= 16'b0000001111000000;
		15'h2338: char_row_bitmap <= 16'b0000001111000000;
		15'h2339: char_row_bitmap <= 16'b0000001111000000;
		15'h233a: char_row_bitmap <= 16'b0000001111000000;
		15'h233b: char_row_bitmap <= 16'b0000001111000000;
		15'h233c: char_row_bitmap <= 16'b0000000000000000;
		15'h233d: char_row_bitmap <= 16'b0000000000000000;
		15'h233e: char_row_bitmap <= 16'b0000000000000000;
		15'h233f: char_row_bitmap <= 16'b0000000000000000;
		15'h2340: char_row_bitmap <= 16'b0000000000000000;
		15'h2341: char_row_bitmap <= 16'b0000000000000000;
		15'h2342: char_row_bitmap <= 16'b0000000000000000;
		15'h2343: char_row_bitmap <= 16'b0000000000000000;
		15'h2344: char_row_bitmap <= 16'b0000000111111111;
		15'h2345: char_row_bitmap <= 16'b0000000111111111;
		15'h2346: char_row_bitmap <= 16'b0000000111111111;
		15'h2347: char_row_bitmap <= 16'b0000000111111111;
		15'h2348: char_row_bitmap <= 16'b0000000110000000;
		15'h2349: char_row_bitmap <= 16'b0000000110000000;
		15'h234a: char_row_bitmap <= 16'b0000000110000000;
		15'h234b: char_row_bitmap <= 16'b0000000110000000;
		15'h234c: char_row_bitmap <= 16'b0000000110000000;
		15'h234d: char_row_bitmap <= 16'b0000000110000000;
		15'h234e: char_row_bitmap <= 16'b0000000110000000;
		15'h234f: char_row_bitmap <= 16'b0000000110000000;
		15'h2350: char_row_bitmap <= 16'b0000001111000000;
		15'h2351: char_row_bitmap <= 16'b0000001111000000;
		15'h2352: char_row_bitmap <= 16'b0000001111000000;
		15'h2353: char_row_bitmap <= 16'b0000001111000000;
		15'h2354: char_row_bitmap <= 16'b0000001111000000;
		15'h2355: char_row_bitmap <= 16'b0000001111000000;
		15'h2356: char_row_bitmap <= 16'b0000001111000000;
		15'h2357: char_row_bitmap <= 16'b0000001111000000;
		15'h2358: char_row_bitmap <= 16'b0000001111000000;
		15'h2359: char_row_bitmap <= 16'b1111111111000000;
		15'h235a: char_row_bitmap <= 16'b1111111111000000;
		15'h235b: char_row_bitmap <= 16'b0000000000000000;
		15'h235c: char_row_bitmap <= 16'b0000000000000000;
		15'h235d: char_row_bitmap <= 16'b0000000000000000;
		15'h235e: char_row_bitmap <= 16'b0000000000000000;
		15'h235f: char_row_bitmap <= 16'b0000000000000000;
		15'h2360: char_row_bitmap <= 16'b0000000000000000;
		15'h2361: char_row_bitmap <= 16'b0000000000000000;
		15'h2362: char_row_bitmap <= 16'b0000000000000000;
		15'h2363: char_row_bitmap <= 16'b0000000000000000;
		15'h2364: char_row_bitmap <= 16'b0000000110000000;
		15'h2365: char_row_bitmap <= 16'b0000000110000000;
		15'h2366: char_row_bitmap <= 16'b0000000110000000;
		15'h2367: char_row_bitmap <= 16'b0000000110000000;
		15'h2368: char_row_bitmap <= 16'b0000000110000000;
		15'h2369: char_row_bitmap <= 16'b0000000110000000;
		15'h236a: char_row_bitmap <= 16'b0000000110000000;
		15'h236b: char_row_bitmap <= 16'b0000000110000000;
		15'h236c: char_row_bitmap <= 16'b1111111110000000;
		15'h236d: char_row_bitmap <= 16'b1111111110000000;
		15'h236e: char_row_bitmap <= 16'b1111111110000000;
		15'h236f: char_row_bitmap <= 16'b1111111110000000;
		15'h2370: char_row_bitmap <= 16'b0000000000000000;
		15'h2371: char_row_bitmap <= 16'b0000000000000000;
		15'h2372: char_row_bitmap <= 16'b0000000000000000;
		15'h2373: char_row_bitmap <= 16'b0000000000000000;
		15'h2374: char_row_bitmap <= 16'b0000000000000000;
		15'h2375: char_row_bitmap <= 16'b0000000000000000;
		15'h2376: char_row_bitmap <= 16'b0000000000000000;
		15'h2377: char_row_bitmap <= 16'b0000000000000000;
		15'h2378: char_row_bitmap <= 16'b0000000000000000;
		15'h2379: char_row_bitmap <= 16'b0000000000000000;
		15'h237a: char_row_bitmap <= 16'b0000000000000000;
		15'h237b: char_row_bitmap <= 16'b0000000000000000;
		15'h237c: char_row_bitmap <= 16'b0000000000000000;
		15'h237d: char_row_bitmap <= 16'b0000000000000000;
		15'h237e: char_row_bitmap <= 16'b0000000000000000;
		15'h237f: char_row_bitmap <= 16'b0000000000000000;
		15'h2380: char_row_bitmap <= 16'b0000000000000000;
		15'h2381: char_row_bitmap <= 16'b1111111111000000;
		15'h2382: char_row_bitmap <= 16'b1111111111000000;
		15'h2383: char_row_bitmap <= 16'b0000001111000000;
		15'h2384: char_row_bitmap <= 16'b0000001111000000;
		15'h2385: char_row_bitmap <= 16'b0000001111000000;
		15'h2386: char_row_bitmap <= 16'b0000001111000000;
		15'h2387: char_row_bitmap <= 16'b0000001111000000;
		15'h2388: char_row_bitmap <= 16'b0000001111000000;
		15'h2389: char_row_bitmap <= 16'b0000001111000000;
		15'h238a: char_row_bitmap <= 16'b0000001111000000;
		15'h238b: char_row_bitmap <= 16'b0000001111000000;
		15'h238c: char_row_bitmap <= 16'b0000000000000000;
		15'h238d: char_row_bitmap <= 16'b0000000000000000;
		15'h238e: char_row_bitmap <= 16'b0000000000000000;
		15'h238f: char_row_bitmap <= 16'b0000000000000000;
		15'h2390: char_row_bitmap <= 16'b0000000000000000;
		15'h2391: char_row_bitmap <= 16'b0000000000000000;
		15'h2392: char_row_bitmap <= 16'b0000000000000000;
		15'h2393: char_row_bitmap <= 16'b0000000000000000;
		15'h2394: char_row_bitmap <= 16'b1111111110000000;
		15'h2395: char_row_bitmap <= 16'b1111111110000000;
		15'h2396: char_row_bitmap <= 16'b1111111110000000;
		15'h2397: char_row_bitmap <= 16'b1111111110000000;
		15'h2398: char_row_bitmap <= 16'b0000000110000000;
		15'h2399: char_row_bitmap <= 16'b0000000110000000;
		15'h239a: char_row_bitmap <= 16'b0000000110000000;
		15'h239b: char_row_bitmap <= 16'b0000000110000000;
		15'h239c: char_row_bitmap <= 16'b0000000110000000;
		15'h239d: char_row_bitmap <= 16'b0000000110000000;
		15'h239e: char_row_bitmap <= 16'b0000000110000000;
		15'h239f: char_row_bitmap <= 16'b0000000110000000;
		15'h23a0: char_row_bitmap <= 16'b0000001111000000;
		15'h23a1: char_row_bitmap <= 16'b0000001111000000;
		15'h23a2: char_row_bitmap <= 16'b0000001111000000;
		15'h23a3: char_row_bitmap <= 16'b0000001111000000;
		15'h23a4: char_row_bitmap <= 16'b0000001111000000;
		15'h23a5: char_row_bitmap <= 16'b0000001111000000;
		15'h23a6: char_row_bitmap <= 16'b0000001111000000;
		15'h23a7: char_row_bitmap <= 16'b0000001111000000;
		15'h23a8: char_row_bitmap <= 16'b0000001111000000;
		15'h23a9: char_row_bitmap <= 16'b0000001111111111;
		15'h23aa: char_row_bitmap <= 16'b0000001111111111;
		15'h23ab: char_row_bitmap <= 16'b0000001111000000;
		15'h23ac: char_row_bitmap <= 16'b0000001111000000;
		15'h23ad: char_row_bitmap <= 16'b0000001111000000;
		15'h23ae: char_row_bitmap <= 16'b0000001111000000;
		15'h23af: char_row_bitmap <= 16'b0000001111000000;
		15'h23b0: char_row_bitmap <= 16'b0000001111000000;
		15'h23b1: char_row_bitmap <= 16'b0000001111000000;
		15'h23b2: char_row_bitmap <= 16'b0000001111000000;
		15'h23b3: char_row_bitmap <= 16'b0000001111000000;
		15'h23b4: char_row_bitmap <= 16'b0000000110000000;
		15'h23b5: char_row_bitmap <= 16'b0000000110000000;
		15'h23b6: char_row_bitmap <= 16'b0000000110000000;
		15'h23b7: char_row_bitmap <= 16'b0000000110000000;
		15'h23b8: char_row_bitmap <= 16'b0000000110000000;
		15'h23b9: char_row_bitmap <= 16'b0000000110000000;
		15'h23ba: char_row_bitmap <= 16'b0000000110000000;
		15'h23bb: char_row_bitmap <= 16'b0000000110000000;
		15'h23bc: char_row_bitmap <= 16'b0000000111111111;
		15'h23bd: char_row_bitmap <= 16'b0000000111111111;
		15'h23be: char_row_bitmap <= 16'b0000000111111111;
		15'h23bf: char_row_bitmap <= 16'b0000000111111111;
		15'h23c0: char_row_bitmap <= 16'b0000000110000000;
		15'h23c1: char_row_bitmap <= 16'b0000000110000000;
		15'h23c2: char_row_bitmap <= 16'b0000000110000000;
		15'h23c3: char_row_bitmap <= 16'b0000000110000000;
		15'h23c4: char_row_bitmap <= 16'b0000000110000000;
		15'h23c5: char_row_bitmap <= 16'b0000000110000000;
		15'h23c6: char_row_bitmap <= 16'b0000000110000000;
		15'h23c7: char_row_bitmap <= 16'b0000000110000000;
		15'h23c8: char_row_bitmap <= 16'b0000001111000000;
		15'h23c9: char_row_bitmap <= 16'b0000001111000000;
		15'h23ca: char_row_bitmap <= 16'b0000001111000000;
		15'h23cb: char_row_bitmap <= 16'b0000001111000000;
		15'h23cc: char_row_bitmap <= 16'b0000001111000000;
		15'h23cd: char_row_bitmap <= 16'b0000001111000000;
		15'h23ce: char_row_bitmap <= 16'b0000001111000000;
		15'h23cf: char_row_bitmap <= 16'b0000001111000000;
		15'h23d0: char_row_bitmap <= 16'b0000001111000000;
		15'h23d1: char_row_bitmap <= 16'b1111111111000000;
		15'h23d2: char_row_bitmap <= 16'b1111111111000000;
		15'h23d3: char_row_bitmap <= 16'b0000001111000000;
		15'h23d4: char_row_bitmap <= 16'b0000001111000000;
		15'h23d5: char_row_bitmap <= 16'b0000001111000000;
		15'h23d6: char_row_bitmap <= 16'b0000001111000000;
		15'h23d7: char_row_bitmap <= 16'b0000001111000000;
		15'h23d8: char_row_bitmap <= 16'b0000001111000000;
		15'h23d9: char_row_bitmap <= 16'b0000001111000000;
		15'h23da: char_row_bitmap <= 16'b0000001111000000;
		15'h23db: char_row_bitmap <= 16'b0000001111000000;
		15'h23dc: char_row_bitmap <= 16'b0000000110000000;
		15'h23dd: char_row_bitmap <= 16'b0000000110000000;
		15'h23de: char_row_bitmap <= 16'b0000000110000000;
		15'h23df: char_row_bitmap <= 16'b0000000110000000;
		15'h23e0: char_row_bitmap <= 16'b0000000110000000;
		15'h23e1: char_row_bitmap <= 16'b0000000110000000;
		15'h23e2: char_row_bitmap <= 16'b0000000110000000;
		15'h23e3: char_row_bitmap <= 16'b0000000110000000;
		15'h23e4: char_row_bitmap <= 16'b1111111110000000;
		15'h23e5: char_row_bitmap <= 16'b1111111110000000;
		15'h23e6: char_row_bitmap <= 16'b1111111110000000;
		15'h23e7: char_row_bitmap <= 16'b1111111110000000;
		15'h23e8: char_row_bitmap <= 16'b0000000110000000;
		15'h23e9: char_row_bitmap <= 16'b0000000110000000;
		15'h23ea: char_row_bitmap <= 16'b0000000110000000;
		15'h23eb: char_row_bitmap <= 16'b0000000110000000;
		15'h23ec: char_row_bitmap <= 16'b0000000110000000;
		15'h23ed: char_row_bitmap <= 16'b0000000110000000;
		15'h23ee: char_row_bitmap <= 16'b0000000110000000;
		15'h23ef: char_row_bitmap <= 16'b0000000110000000;
		15'h23f0: char_row_bitmap <= 16'b0000000110000000;
		15'h23f1: char_row_bitmap <= 16'b0000000110000000;
		15'h23f2: char_row_bitmap <= 16'b0000000110000000;
		15'h23f3: char_row_bitmap <= 16'b0000000110000000;
		15'h23f4: char_row_bitmap <= 16'b0000000110000000;
		15'h23f5: char_row_bitmap <= 16'b0000000110000000;
		15'h23f6: char_row_bitmap <= 16'b0000000110000000;
		15'h23f7: char_row_bitmap <= 16'b0000000110000000;
		15'h23f8: char_row_bitmap <= 16'b1111111111111111;
		15'h23f9: char_row_bitmap <= 16'b1111111111111111;
		15'h23fa: char_row_bitmap <= 16'b1111111111111111;
		15'h23fb: char_row_bitmap <= 16'b1111111111111111;
		15'h23fc: char_row_bitmap <= 16'b0000000000000000;
		15'h23fd: char_row_bitmap <= 16'b0000000000000000;
		15'h23fe: char_row_bitmap <= 16'b0000000000000000;
		15'h23ff: char_row_bitmap <= 16'b0000000000000000;
		15'h2400: char_row_bitmap <= 16'b0000000000000000;
		15'h2401: char_row_bitmap <= 16'b0000000000000000;
		15'h2402: char_row_bitmap <= 16'b0000000000000000;
		15'h2403: char_row_bitmap <= 16'b0000000000000000;
		15'h2404: char_row_bitmap <= 16'b0000001111000000;
		15'h2405: char_row_bitmap <= 16'b0000001111000000;
		15'h2406: char_row_bitmap <= 16'b0000001111000000;
		15'h2407: char_row_bitmap <= 16'b0000001111000000;
		15'h2408: char_row_bitmap <= 16'b0000001111000000;
		15'h2409: char_row_bitmap <= 16'b0000001111000000;
		15'h240a: char_row_bitmap <= 16'b0000001111000000;
		15'h240b: char_row_bitmap <= 16'b0000001111000000;
		15'h240c: char_row_bitmap <= 16'b0000001111000000;
		15'h240d: char_row_bitmap <= 16'b1111111111111111;
		15'h240e: char_row_bitmap <= 16'b1111111111111111;
		15'h240f: char_row_bitmap <= 16'b0000000000000000;
		15'h2410: char_row_bitmap <= 16'b0000000000000000;
		15'h2411: char_row_bitmap <= 16'b0000000000000000;
		15'h2412: char_row_bitmap <= 16'b0000000000000000;
		15'h2413: char_row_bitmap <= 16'b0000000000000000;
		15'h2414: char_row_bitmap <= 16'b0000000000000000;
		15'h2415: char_row_bitmap <= 16'b0000000000000000;
		15'h2416: char_row_bitmap <= 16'b0000000000000000;
		15'h2417: char_row_bitmap <= 16'b0000000000000000;
		15'h2418: char_row_bitmap <= 16'b0000000000000000;
		15'h2419: char_row_bitmap <= 16'b0000000000000000;
		15'h241a: char_row_bitmap <= 16'b0000000000000000;
		15'h241b: char_row_bitmap <= 16'b0000000000000000;
		15'h241c: char_row_bitmap <= 16'b0000000000000000;
		15'h241d: char_row_bitmap <= 16'b0000000000000000;
		15'h241e: char_row_bitmap <= 16'b0000000000000000;
		15'h241f: char_row_bitmap <= 16'b0000000000000000;
		15'h2420: char_row_bitmap <= 16'b1111111111111111;
		15'h2421: char_row_bitmap <= 16'b1111111111111111;
		15'h2422: char_row_bitmap <= 16'b1111111111111111;
		15'h2423: char_row_bitmap <= 16'b1111111111111111;
		15'h2424: char_row_bitmap <= 16'b0000000110000000;
		15'h2425: char_row_bitmap <= 16'b0000000110000000;
		15'h2426: char_row_bitmap <= 16'b0000000110000000;
		15'h2427: char_row_bitmap <= 16'b0000000110000000;
		15'h2428: char_row_bitmap <= 16'b0000000110000000;
		15'h2429: char_row_bitmap <= 16'b0000000110000000;
		15'h242a: char_row_bitmap <= 16'b0000000110000000;
		15'h242b: char_row_bitmap <= 16'b0000000110000000;
		15'h242c: char_row_bitmap <= 16'b0000000000000000;
		15'h242d: char_row_bitmap <= 16'b0000000000000000;
		15'h242e: char_row_bitmap <= 16'b0000000000000000;
		15'h242f: char_row_bitmap <= 16'b0000000000000000;
		15'h2430: char_row_bitmap <= 16'b0000000000000000;
		15'h2431: char_row_bitmap <= 16'b0000000000000000;
		15'h2432: char_row_bitmap <= 16'b0000000000000000;
		15'h2433: char_row_bitmap <= 16'b0000000000000000;
		15'h2434: char_row_bitmap <= 16'b0000000000000000;
		15'h2435: char_row_bitmap <= 16'b1111111111111111;
		15'h2436: char_row_bitmap <= 16'b1111111111111111;
		15'h2437: char_row_bitmap <= 16'b0000001111000000;
		15'h2438: char_row_bitmap <= 16'b0000001111000000;
		15'h2439: char_row_bitmap <= 16'b0000001111000000;
		15'h243a: char_row_bitmap <= 16'b0000001111000000;
		15'h243b: char_row_bitmap <= 16'b0000001111000000;
		15'h243c: char_row_bitmap <= 16'b0000001111000000;
		15'h243d: char_row_bitmap <= 16'b0000001111000000;
		15'h243e: char_row_bitmap <= 16'b0000001111000000;
		15'h243f: char_row_bitmap <= 16'b0000001111000000;
		15'h2440: char_row_bitmap <= 16'b0000001111000000;
		15'h2441: char_row_bitmap <= 16'b0000001111000000;
		15'h2442: char_row_bitmap <= 16'b0000001111000000;
		15'h2443: char_row_bitmap <= 16'b0000001111000000;
		15'h2444: char_row_bitmap <= 16'b0000001111000000;
		15'h2445: char_row_bitmap <= 16'b0000001111000000;
		15'h2446: char_row_bitmap <= 16'b0000001111000000;
		15'h2447: char_row_bitmap <= 16'b0000001111000000;
		15'h2448: char_row_bitmap <= 16'b0000001111111111;
		15'h2449: char_row_bitmap <= 16'b0000001111000000;
		15'h244a: char_row_bitmap <= 16'b0000001111000000;
		15'h244b: char_row_bitmap <= 16'b0000001111111111;
		15'h244c: char_row_bitmap <= 16'b0000000000000000;
		15'h244d: char_row_bitmap <= 16'b0000000000000000;
		15'h244e: char_row_bitmap <= 16'b0000000000000000;
		15'h244f: char_row_bitmap <= 16'b0000000000000000;
		15'h2450: char_row_bitmap <= 16'b0000000000000000;
		15'h2451: char_row_bitmap <= 16'b0000000000000000;
		15'h2452: char_row_bitmap <= 16'b0000000000000000;
		15'h2453: char_row_bitmap <= 16'b0000000000000000;
		15'h2454: char_row_bitmap <= 16'b0000001001000000;
		15'h2455: char_row_bitmap <= 16'b0000001001000000;
		15'h2456: char_row_bitmap <= 16'b0000001001000000;
		15'h2457: char_row_bitmap <= 16'b0000001001000000;
		15'h2458: char_row_bitmap <= 16'b0000001001000000;
		15'h2459: char_row_bitmap <= 16'b0000001001000000;
		15'h245a: char_row_bitmap <= 16'b0000001001000000;
		15'h245b: char_row_bitmap <= 16'b0000001001000000;
		15'h245c: char_row_bitmap <= 16'b0000001111111111;
		15'h245d: char_row_bitmap <= 16'b0000001111111111;
		15'h245e: char_row_bitmap <= 16'b0000001111111111;
		15'h245f: char_row_bitmap <= 16'b0000001111111111;
		15'h2460: char_row_bitmap <= 16'b0000000000000000;
		15'h2461: char_row_bitmap <= 16'b0000000000000000;
		15'h2462: char_row_bitmap <= 16'b0000000000000000;
		15'h2463: char_row_bitmap <= 16'b0000000000000000;
		15'h2464: char_row_bitmap <= 16'b0000000000000000;
		15'h2465: char_row_bitmap <= 16'b0000000000000000;
		15'h2466: char_row_bitmap <= 16'b0000000000000000;
		15'h2467: char_row_bitmap <= 16'b0000000000000000;
		15'h2468: char_row_bitmap <= 16'b0000000000000000;
		15'h2469: char_row_bitmap <= 16'b0000000000000000;
		15'h246a: char_row_bitmap <= 16'b0000000000000000;
		15'h246b: char_row_bitmap <= 16'b0000000000000000;
		15'h246c: char_row_bitmap <= 16'b0000000000000000;
		15'h246d: char_row_bitmap <= 16'b0000000000000000;
		15'h246e: char_row_bitmap <= 16'b0000000000000000;
		15'h246f: char_row_bitmap <= 16'b0000000000000000;
		15'h2470: char_row_bitmap <= 16'b0000001111111111;
		15'h2471: char_row_bitmap <= 16'b0000001111000000;
		15'h2472: char_row_bitmap <= 16'b0000001111000000;
		15'h2473: char_row_bitmap <= 16'b0000001111111111;
		15'h2474: char_row_bitmap <= 16'b0000001111000000;
		15'h2475: char_row_bitmap <= 16'b0000001111000000;
		15'h2476: char_row_bitmap <= 16'b0000001111000000;
		15'h2477: char_row_bitmap <= 16'b0000001111000000;
		15'h2478: char_row_bitmap <= 16'b0000001111000000;
		15'h2479: char_row_bitmap <= 16'b0000001111000000;
		15'h247a: char_row_bitmap <= 16'b0000001111000000;
		15'h247b: char_row_bitmap <= 16'b0000001111000000;
		15'h247c: char_row_bitmap <= 16'b0000000000000000;
		15'h247d: char_row_bitmap <= 16'b0000000000000000;
		15'h247e: char_row_bitmap <= 16'b0000000000000000;
		15'h247f: char_row_bitmap <= 16'b0000000000000000;
		15'h2480: char_row_bitmap <= 16'b0000000000000000;
		15'h2481: char_row_bitmap <= 16'b0000000000000000;
		15'h2482: char_row_bitmap <= 16'b0000000000000000;
		15'h2483: char_row_bitmap <= 16'b0000000000000000;
		15'h2484: char_row_bitmap <= 16'b0000001111111111;
		15'h2485: char_row_bitmap <= 16'b0000001111111111;
		15'h2486: char_row_bitmap <= 16'b0000001111111111;
		15'h2487: char_row_bitmap <= 16'b0000001111111111;
		15'h2488: char_row_bitmap <= 16'b0000001001000000;
		15'h2489: char_row_bitmap <= 16'b0000001001000000;
		15'h248a: char_row_bitmap <= 16'b0000001001000000;
		15'h248b: char_row_bitmap <= 16'b0000001001000000;
		15'h248c: char_row_bitmap <= 16'b0000001001000000;
		15'h248d: char_row_bitmap <= 16'b0000001001000000;
		15'h248e: char_row_bitmap <= 16'b0000001001000000;
		15'h248f: char_row_bitmap <= 16'b0000001001000000;
		15'h2490: char_row_bitmap <= 16'b0000001111000000;
		15'h2491: char_row_bitmap <= 16'b0000001111000000;
		15'h2492: char_row_bitmap <= 16'b0000001111000000;
		15'h2493: char_row_bitmap <= 16'b0000001111000000;
		15'h2494: char_row_bitmap <= 16'b0000001111000000;
		15'h2495: char_row_bitmap <= 16'b0000001111000000;
		15'h2496: char_row_bitmap <= 16'b0000001111000000;
		15'h2497: char_row_bitmap <= 16'b0000001111000000;
		15'h2498: char_row_bitmap <= 16'b1111111111000000;
		15'h2499: char_row_bitmap <= 16'b0000001111000000;
		15'h249a: char_row_bitmap <= 16'b0000001111000000;
		15'h249b: char_row_bitmap <= 16'b1111111111000000;
		15'h249c: char_row_bitmap <= 16'b0000000000000000;
		15'h249d: char_row_bitmap <= 16'b0000000000000000;
		15'h249e: char_row_bitmap <= 16'b0000000000000000;
		15'h249f: char_row_bitmap <= 16'b0000000000000000;
		15'h24a0: char_row_bitmap <= 16'b0000000000000000;
		15'h24a1: char_row_bitmap <= 16'b0000000000000000;
		15'h24a2: char_row_bitmap <= 16'b0000000000000000;
		15'h24a3: char_row_bitmap <= 16'b0000000000000000;
		15'h24a4: char_row_bitmap <= 16'b0000001001000000;
		15'h24a5: char_row_bitmap <= 16'b0000001001000000;
		15'h24a6: char_row_bitmap <= 16'b0000001001000000;
		15'h24a7: char_row_bitmap <= 16'b0000001001000000;
		15'h24a8: char_row_bitmap <= 16'b0000001001000000;
		15'h24a9: char_row_bitmap <= 16'b0000001001000000;
		15'h24aa: char_row_bitmap <= 16'b0000001001000000;
		15'h24ab: char_row_bitmap <= 16'b0000001001000000;
		15'h24ac: char_row_bitmap <= 16'b1111111111000000;
		15'h24ad: char_row_bitmap <= 16'b1111111111000000;
		15'h24ae: char_row_bitmap <= 16'b1111111111000000;
		15'h24af: char_row_bitmap <= 16'b1111111111000000;
		15'h24b0: char_row_bitmap <= 16'b0000000000000000;
		15'h24b1: char_row_bitmap <= 16'b0000000000000000;
		15'h24b2: char_row_bitmap <= 16'b0000000000000000;
		15'h24b3: char_row_bitmap <= 16'b0000000000000000;
		15'h24b4: char_row_bitmap <= 16'b0000000000000000;
		15'h24b5: char_row_bitmap <= 16'b0000000000000000;
		15'h24b6: char_row_bitmap <= 16'b0000000000000000;
		15'h24b7: char_row_bitmap <= 16'b0000000000000000;
		15'h24b8: char_row_bitmap <= 16'b0000000000000000;
		15'h24b9: char_row_bitmap <= 16'b0000000000000000;
		15'h24ba: char_row_bitmap <= 16'b0000000000000000;
		15'h24bb: char_row_bitmap <= 16'b0000000000000000;
		15'h24bc: char_row_bitmap <= 16'b0000000000000000;
		15'h24bd: char_row_bitmap <= 16'b0000000000000000;
		15'h24be: char_row_bitmap <= 16'b0000000000000000;
		15'h24bf: char_row_bitmap <= 16'b0000000000000000;
		15'h24c0: char_row_bitmap <= 16'b1111111111000000;
		15'h24c1: char_row_bitmap <= 16'b0000001111000000;
		15'h24c2: char_row_bitmap <= 16'b0000001111000000;
		15'h24c3: char_row_bitmap <= 16'b1111111111000000;
		15'h24c4: char_row_bitmap <= 16'b0000001111000000;
		15'h24c5: char_row_bitmap <= 16'b0000001111000000;
		15'h24c6: char_row_bitmap <= 16'b0000001111000000;
		15'h24c7: char_row_bitmap <= 16'b0000001111000000;
		15'h24c8: char_row_bitmap <= 16'b0000001111000000;
		15'h24c9: char_row_bitmap <= 16'b0000001111000000;
		15'h24ca: char_row_bitmap <= 16'b0000001111000000;
		15'h24cb: char_row_bitmap <= 16'b0000001111000000;
		15'h24cc: char_row_bitmap <= 16'b0000000000000000;
		15'h24cd: char_row_bitmap <= 16'b0000000000000000;
		15'h24ce: char_row_bitmap <= 16'b0000000000000000;
		15'h24cf: char_row_bitmap <= 16'b0000000000000000;
		15'h24d0: char_row_bitmap <= 16'b0000000000000000;
		15'h24d1: char_row_bitmap <= 16'b0000000000000000;
		15'h24d2: char_row_bitmap <= 16'b0000000000000000;
		15'h24d3: char_row_bitmap <= 16'b0000000000000000;
		15'h24d4: char_row_bitmap <= 16'b1111111111000000;
		15'h24d5: char_row_bitmap <= 16'b1111111111000000;
		15'h24d6: char_row_bitmap <= 16'b1111111111000000;
		15'h24d7: char_row_bitmap <= 16'b1111111111000000;
		15'h24d8: char_row_bitmap <= 16'b0000001001000000;
		15'h24d9: char_row_bitmap <= 16'b0000001001000000;
		15'h24da: char_row_bitmap <= 16'b0000001001000000;
		15'h24db: char_row_bitmap <= 16'b0000001001000000;
		15'h24dc: char_row_bitmap <= 16'b0000001001000000;
		15'h24dd: char_row_bitmap <= 16'b0000001001000000;
		15'h24de: char_row_bitmap <= 16'b0000001001000000;
		15'h24df: char_row_bitmap <= 16'b0000001001000000;
		15'h24e0: char_row_bitmap <= 16'b0000001111000000;
		15'h24e1: char_row_bitmap <= 16'b0000001111000000;
		15'h24e2: char_row_bitmap <= 16'b0000001111000000;
		15'h24e3: char_row_bitmap <= 16'b0000001111000000;
		15'h24e4: char_row_bitmap <= 16'b0000001111000000;
		15'h24e5: char_row_bitmap <= 16'b0000001111000000;
		15'h24e6: char_row_bitmap <= 16'b0000001111000000;
		15'h24e7: char_row_bitmap <= 16'b0000001111000000;
		15'h24e8: char_row_bitmap <= 16'b0000001111111111;
		15'h24e9: char_row_bitmap <= 16'b0000001111000000;
		15'h24ea: char_row_bitmap <= 16'b0000001111000000;
		15'h24eb: char_row_bitmap <= 16'b0000001111111111;
		15'h24ec: char_row_bitmap <= 16'b0000001111000000;
		15'h24ed: char_row_bitmap <= 16'b0000001111000000;
		15'h24ee: char_row_bitmap <= 16'b0000001111000000;
		15'h24ef: char_row_bitmap <= 16'b0000001111000000;
		15'h24f0: char_row_bitmap <= 16'b0000001111000000;
		15'h24f1: char_row_bitmap <= 16'b0000001111000000;
		15'h24f2: char_row_bitmap <= 16'b0000001111000000;
		15'h24f3: char_row_bitmap <= 16'b0000001111000000;
		15'h24f4: char_row_bitmap <= 16'b0000001001000000;
		15'h24f5: char_row_bitmap <= 16'b0000001001000000;
		15'h24f6: char_row_bitmap <= 16'b0000001001000000;
		15'h24f7: char_row_bitmap <= 16'b0000001001000000;
		15'h24f8: char_row_bitmap <= 16'b0000001001000000;
		15'h24f9: char_row_bitmap <= 16'b0000001001000000;
		15'h24fa: char_row_bitmap <= 16'b0000001001000000;
		15'h24fb: char_row_bitmap <= 16'b0000001001000000;
		15'h24fc: char_row_bitmap <= 16'b0000001001111111;
		15'h24fd: char_row_bitmap <= 16'b0000001001111111;
		15'h24fe: char_row_bitmap <= 16'b0000001001111111;
		15'h24ff: char_row_bitmap <= 16'b0000001001111111;
		15'h2500: char_row_bitmap <= 16'b0000001001000000;
		15'h2501: char_row_bitmap <= 16'b0000001001000000;
		15'h2502: char_row_bitmap <= 16'b0000001001000000;
		15'h2503: char_row_bitmap <= 16'b0000001001000000;
		15'h2504: char_row_bitmap <= 16'b0000001001000000;
		15'h2505: char_row_bitmap <= 16'b0000001001000000;
		15'h2506: char_row_bitmap <= 16'b0000001001000000;
		15'h2507: char_row_bitmap <= 16'b0000001001000000;
		15'h2508: char_row_bitmap <= 16'b0000001111000000;
		15'h2509: char_row_bitmap <= 16'b0000001111000000;
		15'h250a: char_row_bitmap <= 16'b0000001111000000;
		15'h250b: char_row_bitmap <= 16'b0000001111000000;
		15'h250c: char_row_bitmap <= 16'b0000001111000000;
		15'h250d: char_row_bitmap <= 16'b0000001111000000;
		15'h250e: char_row_bitmap <= 16'b0000001111000000;
		15'h250f: char_row_bitmap <= 16'b0000001111000000;
		15'h2510: char_row_bitmap <= 16'b0000001111111111;
		15'h2511: char_row_bitmap <= 16'b0000001111111111;
		15'h2512: char_row_bitmap <= 16'b0000001111111111;
		15'h2513: char_row_bitmap <= 16'b0000001111111111;
		15'h2514: char_row_bitmap <= 16'b0000001001000000;
		15'h2515: char_row_bitmap <= 16'b0000001001000000;
		15'h2516: char_row_bitmap <= 16'b0000001001000000;
		15'h2517: char_row_bitmap <= 16'b0000001001000000;
		15'h2518: char_row_bitmap <= 16'b0000001001000000;
		15'h2519: char_row_bitmap <= 16'b0000001001000000;
		15'h251a: char_row_bitmap <= 16'b0000001001000000;
		15'h251b: char_row_bitmap <= 16'b0000001001000000;
		15'h251c: char_row_bitmap <= 16'b0000001001000000;
		15'h251d: char_row_bitmap <= 16'b0000001001000000;
		15'h251e: char_row_bitmap <= 16'b0000001001000000;
		15'h251f: char_row_bitmap <= 16'b0000001001000000;
		15'h2520: char_row_bitmap <= 16'b0000001001000000;
		15'h2521: char_row_bitmap <= 16'b0000001001000000;
		15'h2522: char_row_bitmap <= 16'b0000001001000000;
		15'h2523: char_row_bitmap <= 16'b0000001001000000;
		15'h2524: char_row_bitmap <= 16'b0000001111111111;
		15'h2525: char_row_bitmap <= 16'b0000001111111111;
		15'h2526: char_row_bitmap <= 16'b0000001111111111;
		15'h2527: char_row_bitmap <= 16'b0000001111111111;
		15'h2528: char_row_bitmap <= 16'b0000001111000000;
		15'h2529: char_row_bitmap <= 16'b0000001111000000;
		15'h252a: char_row_bitmap <= 16'b0000001111000000;
		15'h252b: char_row_bitmap <= 16'b0000001111000000;
		15'h252c: char_row_bitmap <= 16'b0000001111000000;
		15'h252d: char_row_bitmap <= 16'b0000001111000000;
		15'h252e: char_row_bitmap <= 16'b0000001111000000;
		15'h252f: char_row_bitmap <= 16'b0000001111000000;
		15'h2530: char_row_bitmap <= 16'b0000001111000000;
		15'h2531: char_row_bitmap <= 16'b0000001111000000;
		15'h2532: char_row_bitmap <= 16'b0000001111000000;
		15'h2533: char_row_bitmap <= 16'b0000001111000000;
		15'h2534: char_row_bitmap <= 16'b0000001111000000;
		15'h2535: char_row_bitmap <= 16'b0000001111000000;
		15'h2536: char_row_bitmap <= 16'b0000001111000000;
		15'h2537: char_row_bitmap <= 16'b0000001111000000;
		15'h2538: char_row_bitmap <= 16'b1111111111000000;
		15'h2539: char_row_bitmap <= 16'b0000001111000000;
		15'h253a: char_row_bitmap <= 16'b0000001111000000;
		15'h253b: char_row_bitmap <= 16'b1111111111000000;
		15'h253c: char_row_bitmap <= 16'b0000001111000000;
		15'h253d: char_row_bitmap <= 16'b0000001111000000;
		15'h253e: char_row_bitmap <= 16'b0000001111000000;
		15'h253f: char_row_bitmap <= 16'b0000001111000000;
		15'h2540: char_row_bitmap <= 16'b0000001111000000;
		15'h2541: char_row_bitmap <= 16'b0000001111000000;
		15'h2542: char_row_bitmap <= 16'b0000001111000000;
		15'h2543: char_row_bitmap <= 16'b0000001111000000;
		15'h2544: char_row_bitmap <= 16'b0000001001000000;
		15'h2545: char_row_bitmap <= 16'b0000001001000000;
		15'h2546: char_row_bitmap <= 16'b0000001001000000;
		15'h2547: char_row_bitmap <= 16'b0000001001000000;
		15'h2548: char_row_bitmap <= 16'b0000001001000000;
		15'h2549: char_row_bitmap <= 16'b0000001001000000;
		15'h254a: char_row_bitmap <= 16'b0000001001000000;
		15'h254b: char_row_bitmap <= 16'b0000001001000000;
		15'h254c: char_row_bitmap <= 16'b1111111001000000;
		15'h254d: char_row_bitmap <= 16'b1111111001000000;
		15'h254e: char_row_bitmap <= 16'b1111111001000000;
		15'h254f: char_row_bitmap <= 16'b1111111001000000;
		15'h2550: char_row_bitmap <= 16'b0000001001000000;
		15'h2551: char_row_bitmap <= 16'b0000001001000000;
		15'h2552: char_row_bitmap <= 16'b0000001001000000;
		15'h2553: char_row_bitmap <= 16'b0000001001000000;
		15'h2554: char_row_bitmap <= 16'b0000001001000000;
		15'h2555: char_row_bitmap <= 16'b0000001001000000;
		15'h2556: char_row_bitmap <= 16'b0000001001000000;
		15'h2557: char_row_bitmap <= 16'b0000001001000000;
		15'h2558: char_row_bitmap <= 16'b0000001111000000;
		15'h2559: char_row_bitmap <= 16'b0000001111000000;
		15'h255a: char_row_bitmap <= 16'b0000001111000000;
		15'h255b: char_row_bitmap <= 16'b0000001111000000;
		15'h255c: char_row_bitmap <= 16'b0000001111000000;
		15'h255d: char_row_bitmap <= 16'b0000001111000000;
		15'h255e: char_row_bitmap <= 16'b0000001111000000;
		15'h255f: char_row_bitmap <= 16'b0000001111000000;
		15'h2560: char_row_bitmap <= 16'b1111111111000000;
		15'h2561: char_row_bitmap <= 16'b1111111111000000;
		15'h2562: char_row_bitmap <= 16'b1111111111000000;
		15'h2563: char_row_bitmap <= 16'b1111111111000000;
		15'h2564: char_row_bitmap <= 16'b0000001001000000;
		15'h2565: char_row_bitmap <= 16'b0000001001000000;
		15'h2566: char_row_bitmap <= 16'b0000001001000000;
		15'h2567: char_row_bitmap <= 16'b0000001001000000;
		15'h2568: char_row_bitmap <= 16'b0000001001000000;
		15'h2569: char_row_bitmap <= 16'b0000001001000000;
		15'h256a: char_row_bitmap <= 16'b0000001001000000;
		15'h256b: char_row_bitmap <= 16'b0000001001000000;
		15'h256c: char_row_bitmap <= 16'b0000001001000000;
		15'h256d: char_row_bitmap <= 16'b0000001001000000;
		15'h256e: char_row_bitmap <= 16'b0000001001000000;
		15'h256f: char_row_bitmap <= 16'b0000001001000000;
		15'h2570: char_row_bitmap <= 16'b0000001001000000;
		15'h2571: char_row_bitmap <= 16'b0000001001000000;
		15'h2572: char_row_bitmap <= 16'b0000001001000000;
		15'h2573: char_row_bitmap <= 16'b0000001001000000;
		15'h2574: char_row_bitmap <= 16'b1111111111000000;
		15'h2575: char_row_bitmap <= 16'b1111111111000000;
		15'h2576: char_row_bitmap <= 16'b1111111111000000;
		15'h2577: char_row_bitmap <= 16'b1111111111000000;
		15'h2578: char_row_bitmap <= 16'b0000001111000000;
		15'h2579: char_row_bitmap <= 16'b0000001111000000;
		15'h257a: char_row_bitmap <= 16'b0000001111000000;
		15'h257b: char_row_bitmap <= 16'b0000001111000000;
		15'h257c: char_row_bitmap <= 16'b0000001111000000;
		15'h257d: char_row_bitmap <= 16'b0000001111000000;
		15'h257e: char_row_bitmap <= 16'b0000001111000000;
		15'h257f: char_row_bitmap <= 16'b0000001111000000;
		15'h2580: char_row_bitmap <= 16'b0000001111000000;
		15'h2581: char_row_bitmap <= 16'b0000001111000000;
		15'h2582: char_row_bitmap <= 16'b0000001111000000;
		15'h2583: char_row_bitmap <= 16'b0000001111000000;
		15'h2584: char_row_bitmap <= 16'b0000001111000000;
		15'h2585: char_row_bitmap <= 16'b0000001111000000;
		15'h2586: char_row_bitmap <= 16'b0000001111000000;
		15'h2587: char_row_bitmap <= 16'b0000001111000000;
		15'h2588: char_row_bitmap <= 16'b1111111111111111;
		15'h2589: char_row_bitmap <= 16'b0000001111111111;
		15'h258a: char_row_bitmap <= 16'b0000001111111111;
		15'h258b: char_row_bitmap <= 16'b1111111111111111;
		15'h258c: char_row_bitmap <= 16'b0000001001000000;
		15'h258d: char_row_bitmap <= 16'b0000001001000000;
		15'h258e: char_row_bitmap <= 16'b0000001001000000;
		15'h258f: char_row_bitmap <= 16'b0000001001000000;
		15'h2590: char_row_bitmap <= 16'b0000001001000000;
		15'h2591: char_row_bitmap <= 16'b0000001001000000;
		15'h2592: char_row_bitmap <= 16'b0000001001000000;
		15'h2593: char_row_bitmap <= 16'b0000001001000000;
		15'h2594: char_row_bitmap <= 16'b0000001111000000;
		15'h2595: char_row_bitmap <= 16'b0000001111000000;
		15'h2596: char_row_bitmap <= 16'b0000001111000000;
		15'h2597: char_row_bitmap <= 16'b0000001111000000;
		15'h2598: char_row_bitmap <= 16'b0000001111000000;
		15'h2599: char_row_bitmap <= 16'b0000001111000000;
		15'h259a: char_row_bitmap <= 16'b0000001111000000;
		15'h259b: char_row_bitmap <= 16'b0000001111000000;
		15'h259c: char_row_bitmap <= 16'b1111111111111111;
		15'h259d: char_row_bitmap <= 16'b1111111111000000;
		15'h259e: char_row_bitmap <= 16'b1111111111000000;
		15'h259f: char_row_bitmap <= 16'b1111111111111111;
		15'h25a0: char_row_bitmap <= 16'b0000001001000000;
		15'h25a1: char_row_bitmap <= 16'b0000001001000000;
		15'h25a2: char_row_bitmap <= 16'b0000001001000000;
		15'h25a3: char_row_bitmap <= 16'b0000001001000000;
		15'h25a4: char_row_bitmap <= 16'b0000001001000000;
		15'h25a5: char_row_bitmap <= 16'b0000001001000000;
		15'h25a6: char_row_bitmap <= 16'b0000001001000000;
		15'h25a7: char_row_bitmap <= 16'b0000001001000000;
		15'h25a8: char_row_bitmap <= 16'b0000001001000000;
		15'h25a9: char_row_bitmap <= 16'b0000001001000000;
		15'h25aa: char_row_bitmap <= 16'b0000001001000000;
		15'h25ab: char_row_bitmap <= 16'b0000001001000000;
		15'h25ac: char_row_bitmap <= 16'b0000001001000000;
		15'h25ad: char_row_bitmap <= 16'b0000001001000000;
		15'h25ae: char_row_bitmap <= 16'b0000001001000000;
		15'h25af: char_row_bitmap <= 16'b0000001001000000;
		15'h25b0: char_row_bitmap <= 16'b1111111111111111;
		15'h25b1: char_row_bitmap <= 16'b1111111111111111;
		15'h25b2: char_row_bitmap <= 16'b1111111111111111;
		15'h25b3: char_row_bitmap <= 16'b1111111111111111;
		15'h25b4: char_row_bitmap <= 16'b0000001111000000;
		15'h25b5: char_row_bitmap <= 16'b0000001111000000;
		15'h25b6: char_row_bitmap <= 16'b0000001111000000;
		15'h25b7: char_row_bitmap <= 16'b0000001111000000;
		15'h25b8: char_row_bitmap <= 16'b0000001111000000;
		15'h25b9: char_row_bitmap <= 16'b0000001111000000;
		15'h25ba: char_row_bitmap <= 16'b0000001111000000;
		15'h25bb: char_row_bitmap <= 16'b0000001111000000;
		15'h25bc: char_row_bitmap <= 16'b0000001111000000;
		15'h25bd: char_row_bitmap <= 16'b0000001111000000;
		15'h25be: char_row_bitmap <= 16'b0000001111000000;
		15'h25bf: char_row_bitmap <= 16'b0000001111000000;
		15'h25c0: char_row_bitmap <= 16'b0000001111000000;
		15'h25c1: char_row_bitmap <= 16'b0000001111000000;
		15'h25c2: char_row_bitmap <= 16'b0000001111000000;
		15'h25c3: char_row_bitmap <= 16'b0000001111000000;
		15'h25c4: char_row_bitmap <= 16'b1111111111111111;
		15'h25c5: char_row_bitmap <= 16'b0000001111111111;
		15'h25c6: char_row_bitmap <= 16'b0000001111111111;
		15'h25c7: char_row_bitmap <= 16'b1111111111111111;
		15'h25c8: char_row_bitmap <= 16'b0000001111000000;
		15'h25c9: char_row_bitmap <= 16'b0000001111000000;
		15'h25ca: char_row_bitmap <= 16'b0000001111000000;
		15'h25cb: char_row_bitmap <= 16'b0000001111000000;
		15'h25cc: char_row_bitmap <= 16'b0000001111000000;
		15'h25cd: char_row_bitmap <= 16'b0000001111000000;
		15'h25ce: char_row_bitmap <= 16'b0000001111000000;
		15'h25cf: char_row_bitmap <= 16'b0000001111000000;
		15'h25d0: char_row_bitmap <= 16'b0000001111000000;
		15'h25d1: char_row_bitmap <= 16'b0000001111000000;
		15'h25d2: char_row_bitmap <= 16'b0000001111000000;
		15'h25d3: char_row_bitmap <= 16'b0000001111000000;
		15'h25d4: char_row_bitmap <= 16'b0000001111000000;
		15'h25d5: char_row_bitmap <= 16'b0000001111000000;
		15'h25d6: char_row_bitmap <= 16'b0000001111000000;
		15'h25d7: char_row_bitmap <= 16'b0000001111000000;
		15'h25d8: char_row_bitmap <= 16'b1111111111111111;
		15'h25d9: char_row_bitmap <= 16'b1111111111111111;
		15'h25da: char_row_bitmap <= 16'b1111111111111111;
		15'h25db: char_row_bitmap <= 16'b1111111111111111;
		15'h25dc: char_row_bitmap <= 16'b0000001001000000;
		15'h25dd: char_row_bitmap <= 16'b0000001001000000;
		15'h25de: char_row_bitmap <= 16'b0000001001000000;
		15'h25df: char_row_bitmap <= 16'b0000001001000000;
		15'h25e0: char_row_bitmap <= 16'b0000001001000000;
		15'h25e1: char_row_bitmap <= 16'b0000001001000000;
		15'h25e2: char_row_bitmap <= 16'b0000001001000000;
		15'h25e3: char_row_bitmap <= 16'b0000001001000000;
		15'h25e4: char_row_bitmap <= 16'b0000001111000000;
		15'h25e5: char_row_bitmap <= 16'b0000001111000000;
		15'h25e6: char_row_bitmap <= 16'b0000001111000000;
		15'h25e7: char_row_bitmap <= 16'b0000001111000000;
		15'h25e8: char_row_bitmap <= 16'b0000001111000000;
		15'h25e9: char_row_bitmap <= 16'b0000001111000000;
		15'h25ea: char_row_bitmap <= 16'b0000001111000000;
		15'h25eb: char_row_bitmap <= 16'b0000001111000000;
		15'h25ec: char_row_bitmap <= 16'b1111111111111111;
		15'h25ed: char_row_bitmap <= 16'b1111111111000000;
		15'h25ee: char_row_bitmap <= 16'b1111111111000000;
		15'h25ef: char_row_bitmap <= 16'b1111111111111111;
		15'h25f0: char_row_bitmap <= 16'b0000001111000000;
		15'h25f1: char_row_bitmap <= 16'b0000001111000000;
		15'h25f2: char_row_bitmap <= 16'b0000001111000000;
		15'h25f3: char_row_bitmap <= 16'b0000001111000000;
		15'h25f4: char_row_bitmap <= 16'b0000001111000000;
		15'h25f5: char_row_bitmap <= 16'b0000001111000000;
		15'h25f6: char_row_bitmap <= 16'b0000001111000000;
		15'h25f7: char_row_bitmap <= 16'b0000001111000000;
		15'h25f8: char_row_bitmap <= 16'b0000001111000000;
		15'h25f9: char_row_bitmap <= 16'b0000001111000000;
		15'h25fa: char_row_bitmap <= 16'b0000001111000000;
		15'h25fb: char_row_bitmap <= 16'b0000001111000000;
		15'h25fc: char_row_bitmap <= 16'b0000001111000000;
		15'h25fd: char_row_bitmap <= 16'b0000001111000000;
		15'h25fe: char_row_bitmap <= 16'b0000001111000000;
		15'h25ff: char_row_bitmap <= 16'b0000001111000000;
		15'h2600: char_row_bitmap <= 16'b1111111111111111;
		15'h2601: char_row_bitmap <= 16'b0000000000000000;
		15'h2602: char_row_bitmap <= 16'b0000000000000000;
		15'h2603: char_row_bitmap <= 16'b1111111111111111;
		15'h2604: char_row_bitmap <= 16'b0000001111000000;
		15'h2605: char_row_bitmap <= 16'b0000001111000000;
		15'h2606: char_row_bitmap <= 16'b0000001111000000;
		15'h2607: char_row_bitmap <= 16'b0000001111000000;
		15'h2608: char_row_bitmap <= 16'b0000001111000000;
		15'h2609: char_row_bitmap <= 16'b0000001111000000;
		15'h260a: char_row_bitmap <= 16'b0000001111000000;
		15'h260b: char_row_bitmap <= 16'b0000001111000000;
		15'h260c: char_row_bitmap <= 16'b0000001001000000;
		15'h260d: char_row_bitmap <= 16'b0000001001000000;
		15'h260e: char_row_bitmap <= 16'b0000001001000000;
		15'h260f: char_row_bitmap <= 16'b0000001001000000;
		15'h2610: char_row_bitmap <= 16'b0000001001000000;
		15'h2611: char_row_bitmap <= 16'b0000001001000000;
		15'h2612: char_row_bitmap <= 16'b0000001001000000;
		15'h2613: char_row_bitmap <= 16'b0000001001000000;
		15'h2614: char_row_bitmap <= 16'b1111111001111111;
		15'h2615: char_row_bitmap <= 16'b1111111001111111;
		15'h2616: char_row_bitmap <= 16'b1111111001111111;
		15'h2617: char_row_bitmap <= 16'b1111111001111111;
		15'h2618: char_row_bitmap <= 16'b0000001001000000;
		15'h2619: char_row_bitmap <= 16'b0000001001000000;
		15'h261a: char_row_bitmap <= 16'b0000001001000000;
		15'h261b: char_row_bitmap <= 16'b0000001001000000;
		15'h261c: char_row_bitmap <= 16'b0000001001000000;
		15'h261d: char_row_bitmap <= 16'b0000001001000000;
		15'h261e: char_row_bitmap <= 16'b0000001001000000;
		15'h261f: char_row_bitmap <= 16'b0000001001000000;
		15'h2620: char_row_bitmap <= 16'b0000001111000000;
		15'h2621: char_row_bitmap <= 16'b0000001111000000;
		15'h2622: char_row_bitmap <= 16'b0000001111000000;
		15'h2623: char_row_bitmap <= 16'b0000001111000000;
		15'h2624: char_row_bitmap <= 16'b0000001111000000;
		15'h2625: char_row_bitmap <= 16'b0000001111000000;
		15'h2626: char_row_bitmap <= 16'b0000001111000000;
		15'h2627: char_row_bitmap <= 16'b0000001111000000;
		15'h2628: char_row_bitmap <= 16'b1111111111111111;
		15'h2629: char_row_bitmap <= 16'b0000000000000000;
		15'h262a: char_row_bitmap <= 16'b0000000000000000;
		15'h262b: char_row_bitmap <= 16'b1111111111111111;
		15'h262c: char_row_bitmap <= 16'b0000000000000000;
		15'h262d: char_row_bitmap <= 16'b0000000000000000;
		15'h262e: char_row_bitmap <= 16'b0000000000000000;
		15'h262f: char_row_bitmap <= 16'b0000000000000000;
		15'h2630: char_row_bitmap <= 16'b0000000000000000;
		15'h2631: char_row_bitmap <= 16'b0000000000000000;
		15'h2632: char_row_bitmap <= 16'b0000000000000000;
		15'h2633: char_row_bitmap <= 16'b0000000000000000;
		15'h2634: char_row_bitmap <= 16'b0000001001000000;
		15'h2635: char_row_bitmap <= 16'b0000001001000000;
		15'h2636: char_row_bitmap <= 16'b0000001001000000;
		15'h2637: char_row_bitmap <= 16'b0000001001000000;
		15'h2638: char_row_bitmap <= 16'b0000001001000000;
		15'h2639: char_row_bitmap <= 16'b0000001001000000;
		15'h263a: char_row_bitmap <= 16'b0000001001000000;
		15'h263b: char_row_bitmap <= 16'b0000001001000000;
		15'h263c: char_row_bitmap <= 16'b1111111111111111;
		15'h263d: char_row_bitmap <= 16'b1111111111111111;
		15'h263e: char_row_bitmap <= 16'b1111111111111111;
		15'h263f: char_row_bitmap <= 16'b1111111111111111;
		15'h2640: char_row_bitmap <= 16'b0000000000000000;
		15'h2641: char_row_bitmap <= 16'b0000000000000000;
		15'h2642: char_row_bitmap <= 16'b0000000000000000;
		15'h2643: char_row_bitmap <= 16'b0000000000000000;
		15'h2644: char_row_bitmap <= 16'b0000000000000000;
		15'h2645: char_row_bitmap <= 16'b0000000000000000;
		15'h2646: char_row_bitmap <= 16'b0000000000000000;
		15'h2647: char_row_bitmap <= 16'b0000000000000000;
		15'h2648: char_row_bitmap <= 16'b0000001111000000;
		15'h2649: char_row_bitmap <= 16'b0000001111000000;
		15'h264a: char_row_bitmap <= 16'b0000001111000000;
		15'h264b: char_row_bitmap <= 16'b0000001111000000;
		15'h264c: char_row_bitmap <= 16'b0000001111000000;
		15'h264d: char_row_bitmap <= 16'b0000001111000000;
		15'h264e: char_row_bitmap <= 16'b0000001111000000;
		15'h264f: char_row_bitmap <= 16'b0000001111000000;
		15'h2650: char_row_bitmap <= 16'b1111111111111111;
		15'h2651: char_row_bitmap <= 16'b1111111111000000;
		15'h2652: char_row_bitmap <= 16'b1111111111000000;
		15'h2653: char_row_bitmap <= 16'b1111111111111111;
		15'h2654: char_row_bitmap <= 16'b0000000000000000;
		15'h2655: char_row_bitmap <= 16'b0000000000000000;
		15'h2656: char_row_bitmap <= 16'b0000000000000000;
		15'h2657: char_row_bitmap <= 16'b0000000000000000;
		15'h2658: char_row_bitmap <= 16'b0000000000000000;
		15'h2659: char_row_bitmap <= 16'b0000000000000000;
		15'h265a: char_row_bitmap <= 16'b0000000000000000;
		15'h265b: char_row_bitmap <= 16'b0000000000000000;
		15'h265c: char_row_bitmap <= 16'b0000001111000000;
		15'h265d: char_row_bitmap <= 16'b0000001111000000;
		15'h265e: char_row_bitmap <= 16'b0000001111000000;
		15'h265f: char_row_bitmap <= 16'b0000001111000000;
		15'h2660: char_row_bitmap <= 16'b0000001111000000;
		15'h2661: char_row_bitmap <= 16'b0000001111000000;
		15'h2662: char_row_bitmap <= 16'b0000001111000000;
		15'h2663: char_row_bitmap <= 16'b0000001111000000;
		15'h2664: char_row_bitmap <= 16'b1111111111111111;
		15'h2665: char_row_bitmap <= 16'b0000001111111111;
		15'h2666: char_row_bitmap <= 16'b0000001111111111;
		15'h2667: char_row_bitmap <= 16'b1111111111111111;
		15'h2668: char_row_bitmap <= 16'b0000000000000000;
		15'h2669: char_row_bitmap <= 16'b0000000000000000;
		15'h266a: char_row_bitmap <= 16'b0000000000000000;
		15'h266b: char_row_bitmap <= 16'b0000000000000000;
		15'h266c: char_row_bitmap <= 16'b0000000000000000;
		15'h266d: char_row_bitmap <= 16'b0000000000000000;
		15'h266e: char_row_bitmap <= 16'b0000000000000000;
		15'h266f: char_row_bitmap <= 16'b0000000000000000;
		15'h2670: char_row_bitmap <= 16'b0000000000000000;
		15'h2671: char_row_bitmap <= 16'b0000000000000000;
		15'h2672: char_row_bitmap <= 16'b0000000000000000;
		15'h2673: char_row_bitmap <= 16'b0000000000000000;
		15'h2674: char_row_bitmap <= 16'b0000000000000000;
		15'h2675: char_row_bitmap <= 16'b0000000000000000;
		15'h2676: char_row_bitmap <= 16'b0000000000000000;
		15'h2677: char_row_bitmap <= 16'b0000000000000000;
		15'h2678: char_row_bitmap <= 16'b1111111111111111;
		15'h2679: char_row_bitmap <= 16'b0000001111111111;
		15'h267a: char_row_bitmap <= 16'b0000001111111111;
		15'h267b: char_row_bitmap <= 16'b1111111111111111;
		15'h267c: char_row_bitmap <= 16'b0000001111000000;
		15'h267d: char_row_bitmap <= 16'b0000001111000000;
		15'h267e: char_row_bitmap <= 16'b0000001111000000;
		15'h267f: char_row_bitmap <= 16'b0000001111000000;
		15'h2680: char_row_bitmap <= 16'b0000001111000000;
		15'h2681: char_row_bitmap <= 16'b0000001111000000;
		15'h2682: char_row_bitmap <= 16'b0000001111000000;
		15'h2683: char_row_bitmap <= 16'b0000001111000000;
		15'h2684: char_row_bitmap <= 16'b0000000000000000;
		15'h2685: char_row_bitmap <= 16'b0000000000000000;
		15'h2686: char_row_bitmap <= 16'b0000000000000000;
		15'h2687: char_row_bitmap <= 16'b0000000000000000;
		15'h2688: char_row_bitmap <= 16'b0000000000000000;
		15'h2689: char_row_bitmap <= 16'b0000000000000000;
		15'h268a: char_row_bitmap <= 16'b0000000000000000;
		15'h268b: char_row_bitmap <= 16'b0000000000000000;
		15'h268c: char_row_bitmap <= 16'b1111111111111111;
		15'h268d: char_row_bitmap <= 16'b1111111111000000;
		15'h268e: char_row_bitmap <= 16'b1111111111000000;
		15'h268f: char_row_bitmap <= 16'b1111111111111111;
		15'h2690: char_row_bitmap <= 16'b0000001111000000;
		15'h2691: char_row_bitmap <= 16'b0000001111000000;
		15'h2692: char_row_bitmap <= 16'b0000001111000000;
		15'h2693: char_row_bitmap <= 16'b0000001111000000;
		15'h2694: char_row_bitmap <= 16'b0000001111000000;
		15'h2695: char_row_bitmap <= 16'b0000001111000000;
		15'h2696: char_row_bitmap <= 16'b0000001111000000;
		15'h2697: char_row_bitmap <= 16'b0000001111000000;
		15'h2698: char_row_bitmap <= 16'b0000000000000000;
		15'h2699: char_row_bitmap <= 16'b0000000000000000;
		15'h269a: char_row_bitmap <= 16'b0000000000000000;
		15'h269b: char_row_bitmap <= 16'b0000000000000000;
		15'h269c: char_row_bitmap <= 16'b0000000000000000;
		15'h269d: char_row_bitmap <= 16'b0000000000000000;
		15'h269e: char_row_bitmap <= 16'b0000000000000000;
		15'h269f: char_row_bitmap <= 16'b0000000000000000;
		15'h26a0: char_row_bitmap <= 16'b1111111111111111;
		15'h26a1: char_row_bitmap <= 16'b1111111111111111;
		15'h26a2: char_row_bitmap <= 16'b1111111111111111;
		15'h26a3: char_row_bitmap <= 16'b1111111111111111;
		15'h26a4: char_row_bitmap <= 16'b0000001001000000;
		15'h26a5: char_row_bitmap <= 16'b0000001001000000;
		15'h26a6: char_row_bitmap <= 16'b0000001001000000;
		15'h26a7: char_row_bitmap <= 16'b0000001001000000;
		15'h26a8: char_row_bitmap <= 16'b0000001001000000;
		15'h26a9: char_row_bitmap <= 16'b0000001001000000;
		15'h26aa: char_row_bitmap <= 16'b0000001001000000;
		15'h26ab: char_row_bitmap <= 16'b0000001001000000;
		15'h26ac: char_row_bitmap <= 16'b0000000000000000;
		15'h26ad: char_row_bitmap <= 16'b0000000000000000;
		15'h26ae: char_row_bitmap <= 16'b0000000000000000;
		15'h26af: char_row_bitmap <= 16'b0000000000000000;
		15'h26b0: char_row_bitmap <= 16'b0000000000000000;
		15'h26b1: char_row_bitmap <= 16'b0000000000000000;
		15'h26b2: char_row_bitmap <= 16'b0000000000000000;
		15'h26b3: char_row_bitmap <= 16'b0000000000000000;
		15'h26b4: char_row_bitmap <= 16'b1111111111111111;
		15'h26b5: char_row_bitmap <= 16'b0000000000000000;
		15'h26b6: char_row_bitmap <= 16'b0000000000000000;
		15'h26b7: char_row_bitmap <= 16'b1111111111111111;
		15'h26b8: char_row_bitmap <= 16'b0000001111000000;
		15'h26b9: char_row_bitmap <= 16'b0000001111000000;
		15'h26ba: char_row_bitmap <= 16'b0000001111000000;
		15'h26bb: char_row_bitmap <= 16'b0000001111000000;
		15'h26bc: char_row_bitmap <= 16'b0000001111000000;
		15'h26bd: char_row_bitmap <= 16'b0000001111000000;
		15'h26be: char_row_bitmap <= 16'b0000001111000000;
		15'h26bf: char_row_bitmap <= 16'b0000001111000000;
		15'h26c0: char_row_bitmap <= 16'b0000001001000000;
		15'h26c1: char_row_bitmap <= 16'b0000001001000000;
		15'h26c2: char_row_bitmap <= 16'b0000001001000000;
		15'h26c3: char_row_bitmap <= 16'b0000001001000000;
		15'h26c4: char_row_bitmap <= 16'b0000001001000000;
		15'h26c5: char_row_bitmap <= 16'b0000001001000000;
		15'h26c6: char_row_bitmap <= 16'b0000001001000000;
		15'h26c7: char_row_bitmap <= 16'b0000001001000000;
		15'h26c8: char_row_bitmap <= 16'b1111111111111111;
		15'h26c9: char_row_bitmap <= 16'b1111111111000000;
		15'h26ca: char_row_bitmap <= 16'b1111111111000000;
		15'h26cb: char_row_bitmap <= 16'b1111111111111111;
		15'h26cc: char_row_bitmap <= 16'b0000001111000000;
		15'h26cd: char_row_bitmap <= 16'b0000001111000000;
		15'h26ce: char_row_bitmap <= 16'b0000001111000000;
		15'h26cf: char_row_bitmap <= 16'b0000001111000000;
		15'h26d0: char_row_bitmap <= 16'b0000001111000000;
		15'h26d1: char_row_bitmap <= 16'b0000001111000000;
		15'h26d2: char_row_bitmap <= 16'b0000001111000000;
		15'h26d3: char_row_bitmap <= 16'b0000001111000000;
		15'h26d4: char_row_bitmap <= 16'b0000001001000000;
		15'h26d5: char_row_bitmap <= 16'b0000001001000000;
		15'h26d6: char_row_bitmap <= 16'b0000001001000000;
		15'h26d7: char_row_bitmap <= 16'b0000001001000000;
		15'h26d8: char_row_bitmap <= 16'b0000001001000000;
		15'h26d9: char_row_bitmap <= 16'b0000001001000000;
		15'h26da: char_row_bitmap <= 16'b0000001001000000;
		15'h26db: char_row_bitmap <= 16'b0000001001000000;
		15'h26dc: char_row_bitmap <= 16'b1111111111111111;
		15'h26dd: char_row_bitmap <= 16'b0000001111111111;
		15'h26de: char_row_bitmap <= 16'b0000001111111111;
		15'h26df: char_row_bitmap <= 16'b1111111111111111;
		15'h26e0: char_row_bitmap <= 16'b0000001111000000;
		15'h26e1: char_row_bitmap <= 16'b0000001111000000;
		15'h26e2: char_row_bitmap <= 16'b0000001111000000;
		15'h26e3: char_row_bitmap <= 16'b0000001111000000;
		15'h26e4: char_row_bitmap <= 16'b0000001111000000;
		15'h26e5: char_row_bitmap <= 16'b0000001111000000;
		15'h26e6: char_row_bitmap <= 16'b0000001111000000;
		15'h26e7: char_row_bitmap <= 16'b0000001111000000;
		15'h26e8: char_row_bitmap <= 16'b0000000000000000;
		15'h26e9: char_row_bitmap <= 16'b0000000000000000;
		15'h26ea: char_row_bitmap <= 16'b0000000000000000;
		15'h26eb: char_row_bitmap <= 16'b0000000000000000;
		15'h26ec: char_row_bitmap <= 16'b0000000000000000;
		15'h26ed: char_row_bitmap <= 16'b0000000000000000;
		15'h26ee: char_row_bitmap <= 16'b0000000000000000;
		15'h26ef: char_row_bitmap <= 16'b0000000000000000;
		15'h26f0: char_row_bitmap <= 16'b1111111111111111;
		15'h26f1: char_row_bitmap <= 16'b1111111100000000;
		15'h26f2: char_row_bitmap <= 16'b1111111100000000;
		15'h26f3: char_row_bitmap <= 16'b1111111111111111;
		15'h26f4: char_row_bitmap <= 16'b0000000000000000;
		15'h26f5: char_row_bitmap <= 16'b0000000000000000;
		15'h26f6: char_row_bitmap <= 16'b0000000000000000;
		15'h26f7: char_row_bitmap <= 16'b0000000000000000;
		15'h26f8: char_row_bitmap <= 16'b0000000000000000;
		15'h26f9: char_row_bitmap <= 16'b0000000000000000;
		15'h26fa: char_row_bitmap <= 16'b0000000000000000;
		15'h26fb: char_row_bitmap <= 16'b0000000000000000;
		15'h26fc: char_row_bitmap <= 16'b0000000000000000;
		15'h26fd: char_row_bitmap <= 16'b0000000000000000;
		15'h26fe: char_row_bitmap <= 16'b0000000000000000;
		15'h26ff: char_row_bitmap <= 16'b0000000000000000;
		15'h2700: char_row_bitmap <= 16'b0000000000000000;
		15'h2701: char_row_bitmap <= 16'b0000000000000000;
		15'h2702: char_row_bitmap <= 16'b0000000000000000;
		15'h2703: char_row_bitmap <= 16'b0000000000000000;
		15'h2704: char_row_bitmap <= 16'b1111111111111111;
		15'h2705: char_row_bitmap <= 16'b0000000011111111;
		15'h2706: char_row_bitmap <= 16'b0000000011111111;
		15'h2707: char_row_bitmap <= 16'b1111111111111111;
		15'h2708: char_row_bitmap <= 16'b0000000000000000;
		15'h2709: char_row_bitmap <= 16'b0000000000000000;
		15'h270a: char_row_bitmap <= 16'b0000000000000000;
		15'h270b: char_row_bitmap <= 16'b0000000000000000;
		15'h270c: char_row_bitmap <= 16'b0000000000000000;
		15'h270d: char_row_bitmap <= 16'b0000000000000000;
		15'h270e: char_row_bitmap <= 16'b0000000000000000;
		15'h270f: char_row_bitmap <= 16'b0000000000000000;
		15'h2710: char_row_bitmap <= 16'b0000001001000000;
		15'h2711: char_row_bitmap <= 16'b0000001001000000;
		15'h2712: char_row_bitmap <= 16'b0000001001000000;
		15'h2713: char_row_bitmap <= 16'b0000001001000000;
		15'h2714: char_row_bitmap <= 16'b0000001001000000;
		15'h2715: char_row_bitmap <= 16'b0000001001000000;
		15'h2716: char_row_bitmap <= 16'b0000001001000000;
		15'h2717: char_row_bitmap <= 16'b0000001001000000;
		15'h2718: char_row_bitmap <= 16'b0000001001000000;
		15'h2719: char_row_bitmap <= 16'b0000001001000000;
		15'h271a: char_row_bitmap <= 16'b0000001111000000;
		15'h271b: char_row_bitmap <= 16'b0000001111000000;
		15'h271c: char_row_bitmap <= 16'b0000001111000000;
		15'h271d: char_row_bitmap <= 16'b0000001111000000;
		15'h271e: char_row_bitmap <= 16'b0000001111000000;
		15'h271f: char_row_bitmap <= 16'b0000001111000000;
		15'h2720: char_row_bitmap <= 16'b0000001111000000;
		15'h2721: char_row_bitmap <= 16'b0000001111000000;
		15'h2722: char_row_bitmap <= 16'b0000001111000000;
		15'h2723: char_row_bitmap <= 16'b0000001111000000;
		15'h2724: char_row_bitmap <= 16'b0000001111000000;
		15'h2725: char_row_bitmap <= 16'b0000001111000000;
		15'h2726: char_row_bitmap <= 16'b0000001111000000;
		15'h2727: char_row_bitmap <= 16'b0000001111000000;
		15'h2728: char_row_bitmap <= 16'b0000001111000000;
		15'h2729: char_row_bitmap <= 16'b0000001111000000;
		15'h272a: char_row_bitmap <= 16'b0000001111000000;
		15'h272b: char_row_bitmap <= 16'b0000001111000000;
		15'h272c: char_row_bitmap <= 16'b0000001111000000;
		15'h272d: char_row_bitmap <= 16'b0000001111000000;
		15'h272e: char_row_bitmap <= 16'b0000001001000000;
		15'h272f: char_row_bitmap <= 16'b0000001001000000;
		15'h2730: char_row_bitmap <= 16'b0000001001000000;
		15'h2731: char_row_bitmap <= 16'b0000001001000000;
		15'h2732: char_row_bitmap <= 16'b0000001001000000;
		15'h2733: char_row_bitmap <= 16'b0000001001000000;
		15'h2734: char_row_bitmap <= 16'b0000001001000000;
		15'h2735: char_row_bitmap <= 16'b0000001001000000;
		15'h2736: char_row_bitmap <= 16'b0000001001000000;
		15'h2737: char_row_bitmap <= 16'b0000001001000000;
		15'h2738: char_row_bitmap <= 16'b0000000110000000;
		15'h2739: char_row_bitmap <= 16'b0000000110000000;
		15'h273a: char_row_bitmap <= 16'b0000000110000000;
		15'h273b: char_row_bitmap <= 16'b0000000110000000;
		15'h273c: char_row_bitmap <= 16'b0000000110000000;
		15'h273d: char_row_bitmap <= 16'b0000000110000000;
		15'h273e: char_row_bitmap <= 16'b0000000110000000;
		15'h273f: char_row_bitmap <= 16'b0000000110000000;
		15'h2740: char_row_bitmap <= 16'b0000000111111111;
		15'h2741: char_row_bitmap <= 16'b0000000110000000;
		15'h2742: char_row_bitmap <= 16'b0000000110000000;
		15'h2743: char_row_bitmap <= 16'b0000000111111111;
		15'h2744: char_row_bitmap <= 16'b0000000110000000;
		15'h2745: char_row_bitmap <= 16'b0000000110000000;
		15'h2746: char_row_bitmap <= 16'b0000000110000000;
		15'h2747: char_row_bitmap <= 16'b0000000110000000;
		15'h2748: char_row_bitmap <= 16'b0000000110000000;
		15'h2749: char_row_bitmap <= 16'b0000000110000000;
		15'h274a: char_row_bitmap <= 16'b0000000110000000;
		15'h274b: char_row_bitmap <= 16'b0000000110000000;
		15'h274c: char_row_bitmap <= 16'b0000000110000000;
		15'h274d: char_row_bitmap <= 16'b0000000110000000;
		15'h274e: char_row_bitmap <= 16'b0000000110000000;
		15'h274f: char_row_bitmap <= 16'b0000000110000000;
		15'h2750: char_row_bitmap <= 16'b0000000110000000;
		15'h2751: char_row_bitmap <= 16'b0000000110000000;
		15'h2752: char_row_bitmap <= 16'b0000000110000000;
		15'h2753: char_row_bitmap <= 16'b0000000110000000;
		15'h2754: char_row_bitmap <= 16'b1111111110000000;
		15'h2755: char_row_bitmap <= 16'b0000000110000000;
		15'h2756: char_row_bitmap <= 16'b0000000110000000;
		15'h2757: char_row_bitmap <= 16'b1111111110000000;
		15'h2758: char_row_bitmap <= 16'b0000000110000000;
		15'h2759: char_row_bitmap <= 16'b0000000110000000;
		15'h275a: char_row_bitmap <= 16'b0000000110000000;
		15'h275b: char_row_bitmap <= 16'b0000000110000000;
		15'h275c: char_row_bitmap <= 16'b0000000110000000;
		15'h275d: char_row_bitmap <= 16'b0000000110000000;
		15'h275e: char_row_bitmap <= 16'b0000000110000000;
		15'h275f: char_row_bitmap <= 16'b0000000110000000;
		15'h2760: char_row_bitmap <= 16'b0000001001000000;
		15'h2761: char_row_bitmap <= 16'b0000001001000000;
		15'h2762: char_row_bitmap <= 16'b0000001001000000;
		15'h2763: char_row_bitmap <= 16'b0000001001000000;
		15'h2764: char_row_bitmap <= 16'b0000001001000000;
		15'h2765: char_row_bitmap <= 16'b0000001001000000;
		15'h2766: char_row_bitmap <= 16'b0000001001000000;
		15'h2767: char_row_bitmap <= 16'b0000001001000000;
		15'h2768: char_row_bitmap <= 16'b0000001001000000;
		15'h2769: char_row_bitmap <= 16'b1111111111111111;
		15'h276a: char_row_bitmap <= 16'b1111111111111111;
		15'h276b: char_row_bitmap <= 16'b0000000000000000;
		15'h276c: char_row_bitmap <= 16'b0000000000000000;
		15'h276d: char_row_bitmap <= 16'b0000000000000000;
		15'h276e: char_row_bitmap <= 16'b0000000000000000;
		15'h276f: char_row_bitmap <= 16'b0000000000000000;
		15'h2770: char_row_bitmap <= 16'b0000000000000000;
		15'h2771: char_row_bitmap <= 16'b0000000000000000;
		15'h2772: char_row_bitmap <= 16'b0000000000000000;
		15'h2773: char_row_bitmap <= 16'b0000000000000000;
		15'h2774: char_row_bitmap <= 16'b0000000000000000;
		15'h2775: char_row_bitmap <= 16'b0000000000000000;
		15'h2776: char_row_bitmap <= 16'b0000000000000000;
		15'h2777: char_row_bitmap <= 16'b0000000000000000;
		15'h2778: char_row_bitmap <= 16'b0000000000000000;
		15'h2779: char_row_bitmap <= 16'b0000000000000000;
		15'h277a: char_row_bitmap <= 16'b0000000000000000;
		15'h277b: char_row_bitmap <= 16'b0000000000000000;
		15'h277c: char_row_bitmap <= 16'b0000000000000000;
		15'h277d: char_row_bitmap <= 16'b1111111111111111;
		15'h277e: char_row_bitmap <= 16'b1111111111111111;
		15'h277f: char_row_bitmap <= 16'b0000001001000000;
		15'h2780: char_row_bitmap <= 16'b0000001001000000;
		15'h2781: char_row_bitmap <= 16'b0000001001000000;
		15'h2782: char_row_bitmap <= 16'b0000001001000000;
		15'h2783: char_row_bitmap <= 16'b0000001001000000;
		15'h2784: char_row_bitmap <= 16'b0000001001000000;
		15'h2785: char_row_bitmap <= 16'b0000001001000000;
		15'h2786: char_row_bitmap <= 16'b0000001001000000;
		15'h2787: char_row_bitmap <= 16'b0000001001000000;
		15'h2788: char_row_bitmap <= 16'b0000000000000000;
		15'h2789: char_row_bitmap <= 16'b0000000000000000;
		15'h278a: char_row_bitmap <= 16'b0000000000000000;
		15'h278b: char_row_bitmap <= 16'b0000000000000000;
		15'h278c: char_row_bitmap <= 16'b0000000000000000;
		15'h278d: char_row_bitmap <= 16'b0000000000000000;
		15'h278e: char_row_bitmap <= 16'b0000000000000000;
		15'h278f: char_row_bitmap <= 16'b0000000000000000;
		15'h2790: char_row_bitmap <= 16'b0000001111111111;
		15'h2791: char_row_bitmap <= 16'b0000001000000000;
		15'h2792: char_row_bitmap <= 16'b0000001000000000;
		15'h2793: char_row_bitmap <= 16'b0000001001111111;
		15'h2794: char_row_bitmap <= 16'b0000001001111111;
		15'h2795: char_row_bitmap <= 16'b0000001001111111;
		15'h2796: char_row_bitmap <= 16'b0000001001111111;
		15'h2797: char_row_bitmap <= 16'b0000001001111111;
		15'h2798: char_row_bitmap <= 16'b0000001001111111;
		15'h2799: char_row_bitmap <= 16'b0000001001111111;
		15'h279a: char_row_bitmap <= 16'b0000001001111111;
		15'h279b: char_row_bitmap <= 16'b0000001001111111;
		15'h279c: char_row_bitmap <= 16'b0000001001111111;
		15'h279d: char_row_bitmap <= 16'b0000001001111111;
		15'h279e: char_row_bitmap <= 16'b0000001001111111;
		15'h279f: char_row_bitmap <= 16'b0000001001111111;
		15'h27a0: char_row_bitmap <= 16'b0000001001111111;
		15'h27a1: char_row_bitmap <= 16'b0000001001111111;
		15'h27a2: char_row_bitmap <= 16'b0000001001111111;
		15'h27a3: char_row_bitmap <= 16'b0000001001111111;
		15'h27a4: char_row_bitmap <= 16'b0000001001111111;
		15'h27a5: char_row_bitmap <= 16'b0000001000000000;
		15'h27a6: char_row_bitmap <= 16'b0000001000000000;
		15'h27a7: char_row_bitmap <= 16'b0000001111111111;
		15'h27a8: char_row_bitmap <= 16'b0000000000000000;
		15'h27a9: char_row_bitmap <= 16'b0000000000000000;
		15'h27aa: char_row_bitmap <= 16'b0000000000000000;
		15'h27ab: char_row_bitmap <= 16'b0000000000000000;
		15'h27ac: char_row_bitmap <= 16'b0000000000000000;
		15'h27ad: char_row_bitmap <= 16'b0000000000000000;
		15'h27ae: char_row_bitmap <= 16'b0000000000000000;
		15'h27af: char_row_bitmap <= 16'b0000000000000000;
		15'h27b0: char_row_bitmap <= 16'b1111111001000000;
		15'h27b1: char_row_bitmap <= 16'b1111111001000000;
		15'h27b2: char_row_bitmap <= 16'b1111111001000000;
		15'h27b3: char_row_bitmap <= 16'b1111111001000000;
		15'h27b4: char_row_bitmap <= 16'b1111111001000000;
		15'h27b5: char_row_bitmap <= 16'b1111111001000000;
		15'h27b6: char_row_bitmap <= 16'b1111111001000000;
		15'h27b7: char_row_bitmap <= 16'b1111111001000000;
		15'h27b8: char_row_bitmap <= 16'b1111111001000000;
		15'h27b9: char_row_bitmap <= 16'b0000000001000000;
		15'h27ba: char_row_bitmap <= 16'b0000000001000000;
		15'h27bb: char_row_bitmap <= 16'b1111111111000000;
		15'h27bc: char_row_bitmap <= 16'b0000000000000000;
		15'h27bd: char_row_bitmap <= 16'b0000000000000000;
		15'h27be: char_row_bitmap <= 16'b0000000000000000;
		15'h27bf: char_row_bitmap <= 16'b0000000000000000;
		15'h27c0: char_row_bitmap <= 16'b0000000000000000;
		15'h27c1: char_row_bitmap <= 16'b0000000000000000;
		15'h27c2: char_row_bitmap <= 16'b0000000000000000;
		15'h27c3: char_row_bitmap <= 16'b0000000000000000;
		15'h27c4: char_row_bitmap <= 16'b0000000000000000;
		15'h27c5: char_row_bitmap <= 16'b0000000000000000;
		15'h27c6: char_row_bitmap <= 16'b0000000000000000;
		15'h27c7: char_row_bitmap <= 16'b0000000000000000;
		15'h27c8: char_row_bitmap <= 16'b0000000000000000;
		15'h27c9: char_row_bitmap <= 16'b0000000000000000;
		15'h27ca: char_row_bitmap <= 16'b0000000000000000;
		15'h27cb: char_row_bitmap <= 16'b0000000000000000;
		15'h27cc: char_row_bitmap <= 16'b1111111111000000;
		15'h27cd: char_row_bitmap <= 16'b0000000001000000;
		15'h27ce: char_row_bitmap <= 16'b0000000001000000;
		15'h27cf: char_row_bitmap <= 16'b1111111001000000;
		15'h27d0: char_row_bitmap <= 16'b1111111001000000;
		15'h27d1: char_row_bitmap <= 16'b1111111001000000;
		15'h27d2: char_row_bitmap <= 16'b1111111001000000;
		15'h27d3: char_row_bitmap <= 16'b1111111001000000;
		15'h27d4: char_row_bitmap <= 16'b1111111001000000;
		15'h27d5: char_row_bitmap <= 16'b1111111001000000;
		15'h27d6: char_row_bitmap <= 16'b1111111001000000;
		15'h27d7: char_row_bitmap <= 16'b1111111001000000;
		15'h27d8: char_row_bitmap <= 16'b0000001001111111;
		15'h27d9: char_row_bitmap <= 16'b0000001001111111;
		15'h27da: char_row_bitmap <= 16'b0000001001111111;
		15'h27db: char_row_bitmap <= 16'b0000001001111111;
		15'h27dc: char_row_bitmap <= 16'b0000001001111111;
		15'h27dd: char_row_bitmap <= 16'b0000001001111111;
		15'h27de: char_row_bitmap <= 16'b0000001001111111;
		15'h27df: char_row_bitmap <= 16'b0000001001111111;
		15'h27e0: char_row_bitmap <= 16'b0000001001111111;
		15'h27e1: char_row_bitmap <= 16'b0000001001111111;
		15'h27e2: char_row_bitmap <= 16'b0000001001111111;
		15'h27e3: char_row_bitmap <= 16'b0000001001111111;
		15'h27e4: char_row_bitmap <= 16'b0000001001111111;
		15'h27e5: char_row_bitmap <= 16'b0000001001111111;
		15'h27e6: char_row_bitmap <= 16'b0000001001111111;
		15'h27e7: char_row_bitmap <= 16'b0000001001111111;
		15'h27e8: char_row_bitmap <= 16'b0000001001111111;
		15'h27e9: char_row_bitmap <= 16'b0000001001111111;
		15'h27ea: char_row_bitmap <= 16'b0000001001111111;
		15'h27eb: char_row_bitmap <= 16'b0000001001111111;
		15'h27ec: char_row_bitmap <= 16'b1111111001000000;
		15'h27ed: char_row_bitmap <= 16'b1111111001000000;
		15'h27ee: char_row_bitmap <= 16'b1111111001000000;
		15'h27ef: char_row_bitmap <= 16'b1111111001000000;
		15'h27f0: char_row_bitmap <= 16'b1111111001000000;
		15'h27f1: char_row_bitmap <= 16'b1111111001000000;
		15'h27f2: char_row_bitmap <= 16'b1111111001000000;
		15'h27f3: char_row_bitmap <= 16'b1111111001000000;
		15'h27f4: char_row_bitmap <= 16'b1111111001000000;
		15'h27f5: char_row_bitmap <= 16'b1111111001000000;
		15'h27f6: char_row_bitmap <= 16'b1111111001000000;
		15'h27f7: char_row_bitmap <= 16'b1111111001000000;
		15'h27f8: char_row_bitmap <= 16'b1111111001000000;
		15'h27f9: char_row_bitmap <= 16'b1111111001000000;
		15'h27fa: char_row_bitmap <= 16'b1111111001000000;
		15'h27fb: char_row_bitmap <= 16'b1111111001000000;
		15'h27fc: char_row_bitmap <= 16'b1111111001000000;
		15'h27fd: char_row_bitmap <= 16'b1111111001000000;
		15'h27fe: char_row_bitmap <= 16'b1111111001000000;
		15'h27ff: char_row_bitmap <= 16'b1111111001000000;
		15'h2800: char_row_bitmap <= 16'b0000000000000000;
		15'h2801: char_row_bitmap <= 16'b0000000000000000;
		15'h2802: char_row_bitmap <= 16'b0000000000000000;
		15'h2803: char_row_bitmap <= 16'b0000000000000000;
		15'h2804: char_row_bitmap <= 16'b0000000000000000;
		15'h2805: char_row_bitmap <= 16'b0000000000000000;
		15'h2806: char_row_bitmap <= 16'b0000000000000000;
		15'h2807: char_row_bitmap <= 16'b0000000000000000;
		15'h2808: char_row_bitmap <= 16'b1111111111111111;
		15'h2809: char_row_bitmap <= 16'b0000000000000000;
		15'h280a: char_row_bitmap <= 16'b0000000000000000;
		15'h280b: char_row_bitmap <= 16'b1111111111111111;
		15'h280c: char_row_bitmap <= 16'b1111111111111111;
		15'h280d: char_row_bitmap <= 16'b1111111111111111;
		15'h280e: char_row_bitmap <= 16'b1111111111111111;
		15'h280f: char_row_bitmap <= 16'b1111111111111111;
		15'h2810: char_row_bitmap <= 16'b1111111111111111;
		15'h2811: char_row_bitmap <= 16'b1111111111111111;
		15'h2812: char_row_bitmap <= 16'b1111111111111111;
		15'h2813: char_row_bitmap <= 16'b1111111111111111;
		15'h2814: char_row_bitmap <= 16'b1111111111111111;
		15'h2815: char_row_bitmap <= 16'b1111111111111111;
		15'h2816: char_row_bitmap <= 16'b1111111111111111;
		15'h2817: char_row_bitmap <= 16'b1111111111111111;
		15'h2818: char_row_bitmap <= 16'b1111111111111111;
		15'h2819: char_row_bitmap <= 16'b1111111111111111;
		15'h281a: char_row_bitmap <= 16'b1111111111111111;
		15'h281b: char_row_bitmap <= 16'b1111111111111111;
		15'h281c: char_row_bitmap <= 16'b1111111111111111;
		15'h281d: char_row_bitmap <= 16'b0000000000000000;
		15'h281e: char_row_bitmap <= 16'b0000000000000000;
		15'h281f: char_row_bitmap <= 16'b1111111111111111;
		15'h2820: char_row_bitmap <= 16'b0000000000000000;
		15'h2821: char_row_bitmap <= 16'b0000000000000000;
		15'h2822: char_row_bitmap <= 16'b0000000000000000;
		15'h2823: char_row_bitmap <= 16'b0000000000000000;
		15'h2824: char_row_bitmap <= 16'b0000000000000000;
		15'h2825: char_row_bitmap <= 16'b0000000000000000;
		15'h2826: char_row_bitmap <= 16'b0000000000000000;
		15'h2827: char_row_bitmap <= 16'b0000000000000000;
		15'h2828: char_row_bitmap <= 16'b0000001001111111;
		15'h2829: char_row_bitmap <= 16'b0000001001111111;
		15'h282a: char_row_bitmap <= 16'b0000001001111111;
		15'h282b: char_row_bitmap <= 16'b0000001001111111;
		15'h282c: char_row_bitmap <= 16'b0000001001111111;
		15'h282d: char_row_bitmap <= 16'b0000001001111111;
		15'h282e: char_row_bitmap <= 16'b0000001001111111;
		15'h282f: char_row_bitmap <= 16'b0000001001111111;
		15'h2830: char_row_bitmap <= 16'b0000001001111111;
		15'h2831: char_row_bitmap <= 16'b0000001000000000;
		15'h2832: char_row_bitmap <= 16'b0000001000000000;
		15'h2833: char_row_bitmap <= 16'b0000001001111111;
		15'h2834: char_row_bitmap <= 16'b0000001001000000;
		15'h2835: char_row_bitmap <= 16'b0000001001000000;
		15'h2836: char_row_bitmap <= 16'b0000001001000000;
		15'h2837: char_row_bitmap <= 16'b0000001001000000;
		15'h2838: char_row_bitmap <= 16'b0000001001000000;
		15'h2839: char_row_bitmap <= 16'b0000001001000000;
		15'h283a: char_row_bitmap <= 16'b0000001001000000;
		15'h283b: char_row_bitmap <= 16'b0000001001000000;
		15'h283c: char_row_bitmap <= 16'b1111111001000000;
		15'h283d: char_row_bitmap <= 16'b1111111001000000;
		15'h283e: char_row_bitmap <= 16'b1111111001000000;
		15'h283f: char_row_bitmap <= 16'b1111111001000000;
		15'h2840: char_row_bitmap <= 16'b1111111001000000;
		15'h2841: char_row_bitmap <= 16'b1111111001000000;
		15'h2842: char_row_bitmap <= 16'b1111111001000000;
		15'h2843: char_row_bitmap <= 16'b1111111001000000;
		15'h2844: char_row_bitmap <= 16'b1111111001000000;
		15'h2845: char_row_bitmap <= 16'b0000000001000000;
		15'h2846: char_row_bitmap <= 16'b0000000001000000;
		15'h2847: char_row_bitmap <= 16'b1111111001000000;
		15'h2848: char_row_bitmap <= 16'b0000001001000000;
		15'h2849: char_row_bitmap <= 16'b0000001001000000;
		15'h284a: char_row_bitmap <= 16'b0000001001000000;
		15'h284b: char_row_bitmap <= 16'b0000001001000000;
		15'h284c: char_row_bitmap <= 16'b0000001001000000;
		15'h284d: char_row_bitmap <= 16'b0000001001000000;
		15'h284e: char_row_bitmap <= 16'b0000001001000000;
		15'h284f: char_row_bitmap <= 16'b0000001001000000;
		15'h2850: char_row_bitmap <= 16'b0000000000000000;
		15'h2851: char_row_bitmap <= 16'b0000000000000000;
		15'h2852: char_row_bitmap <= 16'b0000000000000000;
		15'h2853: char_row_bitmap <= 16'b0000000000000000;
		15'h2854: char_row_bitmap <= 16'b0000000000000000;
		15'h2855: char_row_bitmap <= 16'b0000000000000000;
		15'h2856: char_row_bitmap <= 16'b0000000000000000;
		15'h2857: char_row_bitmap <= 16'b0000000000000000;
		15'h2858: char_row_bitmap <= 16'b1111111111111111;
		15'h2859: char_row_bitmap <= 16'b0000000000000000;
		15'h285a: char_row_bitmap <= 16'b0000000000000000;
		15'h285b: char_row_bitmap <= 16'b1111111001111111;
		15'h285c: char_row_bitmap <= 16'b0000001001111111;
		15'h285d: char_row_bitmap <= 16'b0000001001111111;
		15'h285e: char_row_bitmap <= 16'b0000001001111111;
		15'h285f: char_row_bitmap <= 16'b0000001001111111;
		15'h2860: char_row_bitmap <= 16'b0000001001111111;
		15'h2861: char_row_bitmap <= 16'b0000001001111111;
		15'h2862: char_row_bitmap <= 16'b0000001001111111;
		15'h2863: char_row_bitmap <= 16'b0000001001111111;
		15'h2864: char_row_bitmap <= 16'b0000001001111111;
		15'h2865: char_row_bitmap <= 16'b0000001001111111;
		15'h2866: char_row_bitmap <= 16'b0000001001111111;
		15'h2867: char_row_bitmap <= 16'b0000001001111111;
		15'h2868: char_row_bitmap <= 16'b0000001001111111;
		15'h2869: char_row_bitmap <= 16'b0000001001111111;
		15'h286a: char_row_bitmap <= 16'b0000001001111111;
		15'h286b: char_row_bitmap <= 16'b0000001001111111;
		15'h286c: char_row_bitmap <= 16'b1111111001111111;
		15'h286d: char_row_bitmap <= 16'b0000000000000000;
		15'h286e: char_row_bitmap <= 16'b0000000000000000;
		15'h286f: char_row_bitmap <= 16'b1111111111111111;
		15'h2870: char_row_bitmap <= 16'b0000000000000000;
		15'h2871: char_row_bitmap <= 16'b0000000000000000;
		15'h2872: char_row_bitmap <= 16'b0000000000000000;
		15'h2873: char_row_bitmap <= 16'b0000000000000000;
		15'h2874: char_row_bitmap <= 16'b0000000000000000;
		15'h2875: char_row_bitmap <= 16'b0000000000000000;
		15'h2876: char_row_bitmap <= 16'b0000000000000000;
		15'h2877: char_row_bitmap <= 16'b0000000000000000;
		15'h2878: char_row_bitmap <= 16'b0000001001000000;
		15'h2879: char_row_bitmap <= 16'b0000001001000000;
		15'h287a: char_row_bitmap <= 16'b0000001001000000;
		15'h287b: char_row_bitmap <= 16'b0000001001000000;
		15'h287c: char_row_bitmap <= 16'b0000001001000000;
		15'h287d: char_row_bitmap <= 16'b0000001001000000;
		15'h287e: char_row_bitmap <= 16'b0000001001000000;
		15'h287f: char_row_bitmap <= 16'b0000001001000000;
		15'h2880: char_row_bitmap <= 16'b0000001001111111;
		15'h2881: char_row_bitmap <= 16'b0000001000000000;
		15'h2882: char_row_bitmap <= 16'b0000001000000000;
		15'h2883: char_row_bitmap <= 16'b0000001001111111;
		15'h2884: char_row_bitmap <= 16'b0000001001111111;
		15'h2885: char_row_bitmap <= 16'b0000001001111111;
		15'h2886: char_row_bitmap <= 16'b0000001001111111;
		15'h2887: char_row_bitmap <= 16'b0000001001111111;
		15'h2888: char_row_bitmap <= 16'b0000001001111111;
		15'h2889: char_row_bitmap <= 16'b0000001001111111;
		15'h288a: char_row_bitmap <= 16'b0000001001111111;
		15'h288b: char_row_bitmap <= 16'b0000001001111111;
		15'h288c: char_row_bitmap <= 16'b0000001001000000;
		15'h288d: char_row_bitmap <= 16'b0000001001000000;
		15'h288e: char_row_bitmap <= 16'b0000001001000000;
		15'h288f: char_row_bitmap <= 16'b0000001001000000;
		15'h2890: char_row_bitmap <= 16'b0000001001000000;
		15'h2891: char_row_bitmap <= 16'b0000001001000000;
		15'h2892: char_row_bitmap <= 16'b0000001001000000;
		15'h2893: char_row_bitmap <= 16'b0000001001000000;
		15'h2894: char_row_bitmap <= 16'b1111111001000000;
		15'h2895: char_row_bitmap <= 16'b0000000001000000;
		15'h2896: char_row_bitmap <= 16'b0000000001000000;
		15'h2897: char_row_bitmap <= 16'b1111111001000000;
		15'h2898: char_row_bitmap <= 16'b1111111001000000;
		15'h2899: char_row_bitmap <= 16'b1111111001000000;
		15'h289a: char_row_bitmap <= 16'b1111111001000000;
		15'h289b: char_row_bitmap <= 16'b1111111001000000;
		15'h289c: char_row_bitmap <= 16'b1111111001000000;
		15'h289d: char_row_bitmap <= 16'b1111111001000000;
		15'h289e: char_row_bitmap <= 16'b1111111001000000;
		15'h289f: char_row_bitmap <= 16'b1111111001000000;
		15'h28a0: char_row_bitmap <= 16'b0000000000000000;
		15'h28a1: char_row_bitmap <= 16'b0000000000000000;
		15'h28a2: char_row_bitmap <= 16'b0000000000000000;
		15'h28a3: char_row_bitmap <= 16'b0000000000000000;
		15'h28a4: char_row_bitmap <= 16'b0000000000000000;
		15'h28a5: char_row_bitmap <= 16'b0000000000000000;
		15'h28a6: char_row_bitmap <= 16'b0000000000000000;
		15'h28a7: char_row_bitmap <= 16'b0000000000000000;
		15'h28a8: char_row_bitmap <= 16'b1111111111111111;
		15'h28a9: char_row_bitmap <= 16'b0000000000000000;
		15'h28aa: char_row_bitmap <= 16'b0000000000000000;
		15'h28ab: char_row_bitmap <= 16'b1111111001111111;
		15'h28ac: char_row_bitmap <= 16'b1111111001000000;
		15'h28ad: char_row_bitmap <= 16'b1111111001000000;
		15'h28ae: char_row_bitmap <= 16'b1111111001000000;
		15'h28af: char_row_bitmap <= 16'b1111111001000000;
		15'h28b0: char_row_bitmap <= 16'b1111111001000000;
		15'h28b1: char_row_bitmap <= 16'b1111111001000000;
		15'h28b2: char_row_bitmap <= 16'b1111111001000000;
		15'h28b3: char_row_bitmap <= 16'b1111111001000000;
		15'h28b4: char_row_bitmap <= 16'b1111111001000000;
		15'h28b5: char_row_bitmap <= 16'b1111111001000000;
		15'h28b6: char_row_bitmap <= 16'b1111111001000000;
		15'h28b7: char_row_bitmap <= 16'b1111111001000000;
		15'h28b8: char_row_bitmap <= 16'b1111111001000000;
		15'h28b9: char_row_bitmap <= 16'b1111111001000000;
		15'h28ba: char_row_bitmap <= 16'b1111111001000000;
		15'h28bb: char_row_bitmap <= 16'b1111111001000000;
		15'h28bc: char_row_bitmap <= 16'b1111111001111111;
		15'h28bd: char_row_bitmap <= 16'b0000000000000000;
		15'h28be: char_row_bitmap <= 16'b0000000000000000;
		15'h28bf: char_row_bitmap <= 16'b1111111111111111;
		15'h28c0: char_row_bitmap <= 16'b0000000000000000;
		15'h28c1: char_row_bitmap <= 16'b0000000000000000;
		15'h28c2: char_row_bitmap <= 16'b0000000000000000;
		15'h28c3: char_row_bitmap <= 16'b0000000000000000;
		15'h28c4: char_row_bitmap <= 16'b0000000000000000;
		15'h28c5: char_row_bitmap <= 16'b0000000000000000;
		15'h28c6: char_row_bitmap <= 16'b0000000000000000;
		15'h28c7: char_row_bitmap <= 16'b0000000000000000;
		15'h28c8: char_row_bitmap <= 16'b0000000000000000;
		15'h28c9: char_row_bitmap <= 16'b0000000000000000;
		15'h28ca: char_row_bitmap <= 16'b0000000000000000;
		15'h28cb: char_row_bitmap <= 16'b0000000000000000;
		15'h28cc: char_row_bitmap <= 16'b0000000000000000;
		15'h28cd: char_row_bitmap <= 16'b0000000000000000;
		15'h28ce: char_row_bitmap <= 16'b0000000000000000;
		15'h28cf: char_row_bitmap <= 16'b0000000000000000;
		15'h28d0: char_row_bitmap <= 16'b0000000000000000;
		15'h28d1: char_row_bitmap <= 16'b0000000000000000;
		15'h28d2: char_row_bitmap <= 16'b0000000000000000;
		15'h28d3: char_row_bitmap <= 16'b0000000000000000;
		15'h28d4: char_row_bitmap <= 16'b0000000000000000;
		15'h28d5: char_row_bitmap <= 16'b0000000000000000;
		15'h28d6: char_row_bitmap <= 16'b0000000000000000;
		15'h28d7: char_row_bitmap <= 16'b0000000000000000;
		15'h28d8: char_row_bitmap <= 16'b0000000000000000;
		15'h28d9: char_row_bitmap <= 16'b0000000000000000;
		15'h28da: char_row_bitmap <= 16'b0000000000000000;
		15'h28db: char_row_bitmap <= 16'b0000000000000000;
		15'h28dc: char_row_bitmap <= 16'b0000000000000000;
		15'h28dd: char_row_bitmap <= 16'b0000000000000000;
		15'h28de: char_row_bitmap <= 16'b0000000000000000;
		15'h28df: char_row_bitmap <= 16'b0000000000000000;
		15'h28e0: char_row_bitmap <= 16'b0000000000000000;
		15'h28e1: char_row_bitmap <= 16'b0000000000000000;
		15'h28e2: char_row_bitmap <= 16'b0000000000000000;
		15'h28e3: char_row_bitmap <= 16'b0000000000000000;
		15'h28e4: char_row_bitmap <= 16'b0000000000000000;
		15'h28e5: char_row_bitmap <= 16'b0000000000000000;
		15'h28e6: char_row_bitmap <= 16'b0000000000000000;
		15'h28e7: char_row_bitmap <= 16'b0000000000000000;
		15'h28e8: char_row_bitmap <= 16'b0000000000000000;
		15'h28e9: char_row_bitmap <= 16'b0000000000000000;
		15'h28ea: char_row_bitmap <= 16'b0000000000000000;
		15'h28eb: char_row_bitmap <= 16'b0000000000000000;
		15'h28ec: char_row_bitmap <= 16'b0000000000000000;
		15'h28ed: char_row_bitmap <= 16'b0000000000000000;
		15'h28ee: char_row_bitmap <= 16'b0000000000000000;
		15'h28ef: char_row_bitmap <= 16'b0000000000000000;
		15'h28f0: char_row_bitmap <= 16'b0000000000000000;
		15'h28f1: char_row_bitmap <= 16'b0000000000000000;
		15'h28f2: char_row_bitmap <= 16'b0000000000000000;
		15'h28f3: char_row_bitmap <= 16'b0000000000000000;
		15'h28f4: char_row_bitmap <= 16'b0000000000000000;
		15'h28f5: char_row_bitmap <= 16'b0000000000000000;
		15'h28f6: char_row_bitmap <= 16'b0000000000000000;
		15'h28f7: char_row_bitmap <= 16'b0000000000000000;
		15'h28f8: char_row_bitmap <= 16'b0000000000000000;
		15'h28f9: char_row_bitmap <= 16'b0000000000000000;
		15'h28fa: char_row_bitmap <= 16'b0000000000000000;
		15'h28fb: char_row_bitmap <= 16'b0000000000000000;
		15'h28fc: char_row_bitmap <= 16'b0000000000000000;
		15'h28fd: char_row_bitmap <= 16'b0000000000000000;
		15'h28fe: char_row_bitmap <= 16'b0000000000000000;
		15'h28ff: char_row_bitmap <= 16'b0000000000000000;
		15'h2900: char_row_bitmap <= 16'b0000000000000000;
		15'h2901: char_row_bitmap <= 16'b0000000000000000;
		15'h2902: char_row_bitmap <= 16'b0000000000000000;
		15'h2903: char_row_bitmap <= 16'b0000000000000000;
		15'h2904: char_row_bitmap <= 16'b0000000000000000;
		15'h2905: char_row_bitmap <= 16'b0000000000000000;
		15'h2906: char_row_bitmap <= 16'b0000000000000000;
		15'h2907: char_row_bitmap <= 16'b0000000000000000;
		15'h2908: char_row_bitmap <= 16'b0000000000000000;
		15'h2909: char_row_bitmap <= 16'b0000000000000000;
		15'h290a: char_row_bitmap <= 16'b0000000000000000;
		15'h290b: char_row_bitmap <= 16'b0000000000000000;
		15'h290c: char_row_bitmap <= 16'b0000000000000000;
		15'h290d: char_row_bitmap <= 16'b0000000000000000;
		15'h290e: char_row_bitmap <= 16'b0000000000000000;
		15'h290f: char_row_bitmap <= 16'b0000000000000000;
		15'h2910: char_row_bitmap <= 16'b0000000000000000;
		15'h2911: char_row_bitmap <= 16'b0000000000000000;
		15'h2912: char_row_bitmap <= 16'b0000000000000000;
		15'h2913: char_row_bitmap <= 16'b0000000000000000;
		15'h2914: char_row_bitmap <= 16'b0000000000000000;
		15'h2915: char_row_bitmap <= 16'b0000000000000000;
		15'h2916: char_row_bitmap <= 16'b0000000000000000;
		15'h2917: char_row_bitmap <= 16'b0000000000000000;
		15'h2918: char_row_bitmap <= 16'b0000000000000000;
		15'h2919: char_row_bitmap <= 16'b0000000000000000;
		15'h291a: char_row_bitmap <= 16'b0000000000000000;
		15'h291b: char_row_bitmap <= 16'b0000000000000000;
		15'h291c: char_row_bitmap <= 16'b0000000000000000;
		15'h291d: char_row_bitmap <= 16'b0000000000000000;
		15'h291e: char_row_bitmap <= 16'b0000000000000000;
		15'h291f: char_row_bitmap <= 16'b0000000000000000;
		15'h2920: char_row_bitmap <= 16'b0000000000000000;
		15'h2921: char_row_bitmap <= 16'b0000000000000000;
		15'h2922: char_row_bitmap <= 16'b0000000000000000;
		15'h2923: char_row_bitmap <= 16'b0000000000000000;
		15'h2924: char_row_bitmap <= 16'b0000000000000000;
		15'h2925: char_row_bitmap <= 16'b0000000000000000;
		15'h2926: char_row_bitmap <= 16'b0000000000000000;
		15'h2927: char_row_bitmap <= 16'b0000000000000000;
		15'h2928: char_row_bitmap <= 16'b0000000000000000;
		15'h2929: char_row_bitmap <= 16'b0000000000000000;
		15'h292a: char_row_bitmap <= 16'b0000000000000000;
		15'h292b: char_row_bitmap <= 16'b0000000000000000;
		15'h292c: char_row_bitmap <= 16'b0000000000000000;
		15'h292d: char_row_bitmap <= 16'b0000000000000000;
		15'h292e: char_row_bitmap <= 16'b0000000000000000;
		15'h292f: char_row_bitmap <= 16'b0000000000000000;
		15'h2930: char_row_bitmap <= 16'b0000000000000000;
		15'h2931: char_row_bitmap <= 16'b0000000000000000;
		15'h2932: char_row_bitmap <= 16'b0000000000000000;
		15'h2933: char_row_bitmap <= 16'b0000000000000000;
		15'h2934: char_row_bitmap <= 16'b0000000000000000;
		15'h2935: char_row_bitmap <= 16'b0000000000000000;
		15'h2936: char_row_bitmap <= 16'b0000000000000000;
		15'h2937: char_row_bitmap <= 16'b0000000000000000;
		15'h2938: char_row_bitmap <= 16'b0000000000000000;
		15'h2939: char_row_bitmap <= 16'b0000000000000000;
		15'h293a: char_row_bitmap <= 16'b0000000000000000;
		15'h293b: char_row_bitmap <= 16'b0000000000000000;
		15'h293c: char_row_bitmap <= 16'b0000000000000000;
		15'h293d: char_row_bitmap <= 16'b0000000000000000;
		15'h293e: char_row_bitmap <= 16'b0000000000000000;
		15'h293f: char_row_bitmap <= 16'b0000000000000000;
		15'h2940: char_row_bitmap <= 16'b0000000000000000;
		15'h2941: char_row_bitmap <= 16'b0000000011000000;
		15'h2942: char_row_bitmap <= 16'b0000000111100000;
		15'h2943: char_row_bitmap <= 16'b0000001111110000;
		15'h2944: char_row_bitmap <= 16'b0000011111111000;
		15'h2945: char_row_bitmap <= 16'b0000111111111100;
		15'h2946: char_row_bitmap <= 16'b0001111111111110;
		15'h2947: char_row_bitmap <= 16'b0000000111100000;
		15'h2948: char_row_bitmap <= 16'b0000000111100000;
		15'h2949: char_row_bitmap <= 16'b0000001111100000;
		15'h294a: char_row_bitmap <= 16'b0111111111000000;
		15'h294b: char_row_bitmap <= 16'b0111111111000000;
		15'h294c: char_row_bitmap <= 16'b0111111110000000;
		15'h294d: char_row_bitmap <= 16'b0111111000000000;
		15'h294e: char_row_bitmap <= 16'b0000000000000000;
		15'h294f: char_row_bitmap <= 16'b0000000000000000;
		15'h2950: char_row_bitmap <= 16'b0000000000000000;
		15'h2951: char_row_bitmap <= 16'b0000000000000000;
		15'h2952: char_row_bitmap <= 16'b0000000000000000;
		15'h2953: char_row_bitmap <= 16'b0000000000000000;
		15'h2954: char_row_bitmap <= 16'b0000000000000011;
		15'h2955: char_row_bitmap <= 16'b0000000000000111;
		15'h2956: char_row_bitmap <= 16'b0000000000000110;
		15'h2957: char_row_bitmap <= 16'b0000000000001110;
		15'h2958: char_row_bitmap <= 16'b0000000000011100;
		15'h2959: char_row_bitmap <= 16'b0000000000111000;
		15'h295a: char_row_bitmap <= 16'b0000000001110000;
		15'h295b: char_row_bitmap <= 16'b0000000001100000;
		15'h295c: char_row_bitmap <= 16'b0000000011100000;
		15'h295d: char_row_bitmap <= 16'b0000000011000000;
		15'h295e: char_row_bitmap <= 16'b0000000000000000;
		15'h295f: char_row_bitmap <= 16'b0000000000000000;
		15'h2960: char_row_bitmap <= 16'b0000000000000000;
		15'h2961: char_row_bitmap <= 16'b0000000000000000;
		15'h2962: char_row_bitmap <= 16'b0000000000000000;
		15'h2963: char_row_bitmap <= 16'b0000000000000000;
		15'h2964: char_row_bitmap <= 16'b0000000000000000;
		15'h2965: char_row_bitmap <= 16'b0000000000000000;
		15'h2966: char_row_bitmap <= 16'b0000000000000000;
		15'h2967: char_row_bitmap <= 16'b0000000000000000;
		15'h2968: char_row_bitmap <= 16'b0000000000000000;
		15'h2969: char_row_bitmap <= 16'b0000000000000000;
		15'h296a: char_row_bitmap <= 16'b0000000000000000;
		15'h296b: char_row_bitmap <= 16'b0000000000000000;
		15'h296c: char_row_bitmap <= 16'b0000000000000000;
		15'h296d: char_row_bitmap <= 16'b0000000000000000;
		15'h296e: char_row_bitmap <= 16'b0000000000000000;
		15'h296f: char_row_bitmap <= 16'b0000000000000000;
		15'h2970: char_row_bitmap <= 16'b0000000000000000;
		15'h2971: char_row_bitmap <= 16'b0000000000000000;
		15'h2972: char_row_bitmap <= 16'b0000000011000000;
		15'h2973: char_row_bitmap <= 16'b0000000011100000;
		15'h2974: char_row_bitmap <= 16'b0000000001100000;
		15'h2975: char_row_bitmap <= 16'b0000000001110000;
		15'h2976: char_row_bitmap <= 16'b0000000000111000;
		15'h2977: char_row_bitmap <= 16'b0000000000011100;
		15'h2978: char_row_bitmap <= 16'b0000000000001110;
		15'h2979: char_row_bitmap <= 16'b0000000000000110;
		15'h297a: char_row_bitmap <= 16'b0000000000000111;
		15'h297b: char_row_bitmap <= 16'b0000000000000011;
		15'h297c: char_row_bitmap <= 16'b0000000000000000;
		15'h297d: char_row_bitmap <= 16'b0000000000000000;
		15'h297e: char_row_bitmap <= 16'b0000000000000000;
		15'h297f: char_row_bitmap <= 16'b0000000000000000;
		15'h2980: char_row_bitmap <= 16'b0000000000000000;
		15'h2981: char_row_bitmap <= 16'b0000000000000000;
		15'h2982: char_row_bitmap <= 16'b0000000000000000;
		15'h2983: char_row_bitmap <= 16'b0000000000000000;
		15'h2984: char_row_bitmap <= 16'b0000000000000000;
		15'h2985: char_row_bitmap <= 16'b0000000000000000;
		15'h2986: char_row_bitmap <= 16'b0000001100000000;
		15'h2987: char_row_bitmap <= 16'b0000011100000000;
		15'h2988: char_row_bitmap <= 16'b0000011000000000;
		15'h2989: char_row_bitmap <= 16'b0000111000000000;
		15'h298a: char_row_bitmap <= 16'b0001110000000000;
		15'h298b: char_row_bitmap <= 16'b0011100000000000;
		15'h298c: char_row_bitmap <= 16'b0111000000000000;
		15'h298d: char_row_bitmap <= 16'b0110000000000000;
		15'h298e: char_row_bitmap <= 16'b1110000000000000;
		15'h298f: char_row_bitmap <= 16'b1100000000000000;
		15'h2990: char_row_bitmap <= 16'b1100000000000000;
		15'h2991: char_row_bitmap <= 16'b1110000000000000;
		15'h2992: char_row_bitmap <= 16'b0110000000000000;
		15'h2993: char_row_bitmap <= 16'b0111000000000000;
		15'h2994: char_row_bitmap <= 16'b0011100000000000;
		15'h2995: char_row_bitmap <= 16'b0001110000000000;
		15'h2996: char_row_bitmap <= 16'b0000111000000000;
		15'h2997: char_row_bitmap <= 16'b0000011000000000;
		15'h2998: char_row_bitmap <= 16'b0000011100000000;
		15'h2999: char_row_bitmap <= 16'b0000001100000000;
		15'h299a: char_row_bitmap <= 16'b0000000000000000;
		15'h299b: char_row_bitmap <= 16'b0000000000000000;
		15'h299c: char_row_bitmap <= 16'b0000000000000000;
		15'h299d: char_row_bitmap <= 16'b0000000000000000;
		15'h299e: char_row_bitmap <= 16'b0000000000000000;
		15'h299f: char_row_bitmap <= 16'b0000000000000000;
		15'h29a0: char_row_bitmap <= 16'b0000000000000000;
		15'h29a1: char_row_bitmap <= 16'b0000000000000000;
		15'h29a2: char_row_bitmap <= 16'b0000000000000000;
		15'h29a3: char_row_bitmap <= 16'b0000000000000000;
		15'h29a4: char_row_bitmap <= 16'b1100000000000000;
		15'h29a5: char_row_bitmap <= 16'b1110000000000000;
		15'h29a6: char_row_bitmap <= 16'b0110000000000000;
		15'h29a7: char_row_bitmap <= 16'b0011000000000000;
		15'h29a8: char_row_bitmap <= 16'b0011100000000000;
		15'h29a9: char_row_bitmap <= 16'b0001110000000000;
		15'h29aa: char_row_bitmap <= 16'b0000111000000000;
		15'h29ab: char_row_bitmap <= 16'b0000011000000000;
		15'h29ac: char_row_bitmap <= 16'b0000011100000000;
		15'h29ad: char_row_bitmap <= 16'b0000001100000000;
		15'h29ae: char_row_bitmap <= 16'b0000001100000000;
		15'h29af: char_row_bitmap <= 16'b0000011100000000;
		15'h29b0: char_row_bitmap <= 16'b0000011000000000;
		15'h29b1: char_row_bitmap <= 16'b0000111000000000;
		15'h29b2: char_row_bitmap <= 16'b0001110000000000;
		15'h29b3: char_row_bitmap <= 16'b0011100000000000;
		15'h29b4: char_row_bitmap <= 16'b0111000000000000;
		15'h29b5: char_row_bitmap <= 16'b0110000000000000;
		15'h29b6: char_row_bitmap <= 16'b1110000000000000;
		15'h29b7: char_row_bitmap <= 16'b1100000000000000;
		15'h29b8: char_row_bitmap <= 16'b1100000000000011;
		15'h29b9: char_row_bitmap <= 16'b1110000000000111;
		15'h29ba: char_row_bitmap <= 16'b0110000000000110;
		15'h29bb: char_row_bitmap <= 16'b0011000000001100;
		15'h29bc: char_row_bitmap <= 16'b0011100000011100;
		15'h29bd: char_row_bitmap <= 16'b0001110000111000;
		15'h29be: char_row_bitmap <= 16'b0000111001110000;
		15'h29bf: char_row_bitmap <= 16'b0000011001100000;
		15'h29c0: char_row_bitmap <= 16'b0000011111100000;
		15'h29c1: char_row_bitmap <= 16'b0000001111000000;
		15'h29c2: char_row_bitmap <= 16'b0000000000000000;
		15'h29c3: char_row_bitmap <= 16'b0000000000000000;
		15'h29c4: char_row_bitmap <= 16'b0000000000000000;
		15'h29c5: char_row_bitmap <= 16'b0000000000000000;
		15'h29c6: char_row_bitmap <= 16'b0000000000000000;
		15'h29c7: char_row_bitmap <= 16'b0000000000000000;
		15'h29c8: char_row_bitmap <= 16'b0000000000000000;
		15'h29c9: char_row_bitmap <= 16'b0000000000000000;
		15'h29ca: char_row_bitmap <= 16'b0000000000000000;
		15'h29cb: char_row_bitmap <= 16'b0000000000000000;
		15'h29cc: char_row_bitmap <= 16'b0000000000000011;
		15'h29cd: char_row_bitmap <= 16'b0000000000000111;
		15'h29ce: char_row_bitmap <= 16'b0000000000000110;
		15'h29cf: char_row_bitmap <= 16'b0000000000001100;
		15'h29d0: char_row_bitmap <= 16'b0000000000011100;
		15'h29d1: char_row_bitmap <= 16'b0000000000111000;
		15'h29d2: char_row_bitmap <= 16'b0000000001110000;
		15'h29d3: char_row_bitmap <= 16'b0000000001100000;
		15'h29d4: char_row_bitmap <= 16'b0000000011100000;
		15'h29d5: char_row_bitmap <= 16'b0000000011000000;
		15'h29d6: char_row_bitmap <= 16'b0000000011000000;
		15'h29d7: char_row_bitmap <= 16'b0000000011100000;
		15'h29d8: char_row_bitmap <= 16'b0000000001100000;
		15'h29d9: char_row_bitmap <= 16'b0000000001110000;
		15'h29da: char_row_bitmap <= 16'b0000000000111000;
		15'h29db: char_row_bitmap <= 16'b0000000000011100;
		15'h29dc: char_row_bitmap <= 16'b0000000000001110;
		15'h29dd: char_row_bitmap <= 16'b0000000000000110;
		15'h29de: char_row_bitmap <= 16'b0000000000000111;
		15'h29df: char_row_bitmap <= 16'b0000000000000011;
		15'h29e0: char_row_bitmap <= 16'b0000000000000000;
		15'h29e1: char_row_bitmap <= 16'b0000000000000000;
		15'h29e2: char_row_bitmap <= 16'b0000000000000000;
		15'h29e3: char_row_bitmap <= 16'b0000000000000000;
		15'h29e4: char_row_bitmap <= 16'b0000000000000000;
		15'h29e5: char_row_bitmap <= 16'b0000000000000000;
		15'h29e6: char_row_bitmap <= 16'b0000000000000000;
		15'h29e7: char_row_bitmap <= 16'b0000000000000000;
		15'h29e8: char_row_bitmap <= 16'b0000000000000000;
		15'h29e9: char_row_bitmap <= 16'b0000000000000000;
		15'h29ea: char_row_bitmap <= 16'b0000001111000000;
		15'h29eb: char_row_bitmap <= 16'b0000011111100000;
		15'h29ec: char_row_bitmap <= 16'b0000011001100000;
		15'h29ed: char_row_bitmap <= 16'b0000111001110000;
		15'h29ee: char_row_bitmap <= 16'b0001110000111000;
		15'h29ef: char_row_bitmap <= 16'b0011100000011100;
		15'h29f0: char_row_bitmap <= 16'b0111000000001110;
		15'h29f1: char_row_bitmap <= 16'b0110000000000110;
		15'h29f2: char_row_bitmap <= 16'b1110000000000111;
		15'h29f3: char_row_bitmap <= 16'b1100000000000011;
		15'h29f4: char_row_bitmap <= 16'b1100000000000000;
		15'h29f5: char_row_bitmap <= 16'b1110000000000000;
		15'h29f6: char_row_bitmap <= 16'b0110000000000000;
		15'h29f7: char_row_bitmap <= 16'b0011000000000000;
		15'h29f8: char_row_bitmap <= 16'b0011100000000000;
		15'h29f9: char_row_bitmap <= 16'b0001110000000000;
		15'h29fa: char_row_bitmap <= 16'b0000111000000000;
		15'h29fb: char_row_bitmap <= 16'b0000011000000000;
		15'h29fc: char_row_bitmap <= 16'b0000011100000000;
		15'h29fd: char_row_bitmap <= 16'b0000001110000000;
		15'h29fe: char_row_bitmap <= 16'b0000001111000000;
		15'h29ff: char_row_bitmap <= 16'b0000011111100000;
		15'h2a00: char_row_bitmap <= 16'b0000011001100000;
		15'h2a01: char_row_bitmap <= 16'b0000111001110000;
		15'h2a02: char_row_bitmap <= 16'b0001110000111000;
		15'h2a03: char_row_bitmap <= 16'b0011100000011100;
		15'h2a04: char_row_bitmap <= 16'b0111000000001110;
		15'h2a05: char_row_bitmap <= 16'b0110000000000110;
		15'h2a06: char_row_bitmap <= 16'b1110000000000111;
		15'h2a07: char_row_bitmap <= 16'b1100000000000011;
		15'h2a08: char_row_bitmap <= 16'b1100000000000011;
		15'h2a09: char_row_bitmap <= 16'b1110000000000111;
		15'h2a0a: char_row_bitmap <= 16'b0110000000000110;
		15'h2a0b: char_row_bitmap <= 16'b0111000000001110;
		15'h2a0c: char_row_bitmap <= 16'b0011100000011100;
		15'h2a0d: char_row_bitmap <= 16'b0001110000111000;
		15'h2a0e: char_row_bitmap <= 16'b0000111001110000;
		15'h2a0f: char_row_bitmap <= 16'b0000011001100000;
		15'h2a10: char_row_bitmap <= 16'b0000011111100000;
		15'h2a11: char_row_bitmap <= 16'b0000001111000000;
		15'h2a12: char_row_bitmap <= 16'b0000001110000000;
		15'h2a13: char_row_bitmap <= 16'b0000011100000000;
		15'h2a14: char_row_bitmap <= 16'b0000011000000000;
		15'h2a15: char_row_bitmap <= 16'b0000111000000000;
		15'h2a16: char_row_bitmap <= 16'b0001110000000000;
		15'h2a17: char_row_bitmap <= 16'b0011100000000000;
		15'h2a18: char_row_bitmap <= 16'b0011000000000000;
		15'h2a19: char_row_bitmap <= 16'b0110000000000000;
		15'h2a1a: char_row_bitmap <= 16'b1110000000000000;
		15'h2a1b: char_row_bitmap <= 16'b1100000000000000;
		15'h2a1c: char_row_bitmap <= 16'b1100000000000011;
		15'h2a1d: char_row_bitmap <= 16'b1110000000000111;
		15'h2a1e: char_row_bitmap <= 16'b0110000000000110;
		15'h2a1f: char_row_bitmap <= 16'b0111000000001110;
		15'h2a20: char_row_bitmap <= 16'b0011100000011100;
		15'h2a21: char_row_bitmap <= 16'b0001110000111000;
		15'h2a22: char_row_bitmap <= 16'b0000111001110000;
		15'h2a23: char_row_bitmap <= 16'b0000011001100000;
		15'h2a24: char_row_bitmap <= 16'b0000011111100000;
		15'h2a25: char_row_bitmap <= 16'b0000001111000000;
		15'h2a26: char_row_bitmap <= 16'b0000000111000000;
		15'h2a27: char_row_bitmap <= 16'b0000000011100000;
		15'h2a28: char_row_bitmap <= 16'b0000000001100000;
		15'h2a29: char_row_bitmap <= 16'b0000000001110000;
		15'h2a2a: char_row_bitmap <= 16'b0000000000111000;
		15'h2a2b: char_row_bitmap <= 16'b0000000000011100;
		15'h2a2c: char_row_bitmap <= 16'b0000000000001100;
		15'h2a2d: char_row_bitmap <= 16'b0000000000000110;
		15'h2a2e: char_row_bitmap <= 16'b0000000000000111;
		15'h2a2f: char_row_bitmap <= 16'b0000000000000011;
		15'h2a30: char_row_bitmap <= 16'b0000000000000011;
		15'h2a31: char_row_bitmap <= 16'b0000000000000111;
		15'h2a32: char_row_bitmap <= 16'b0000000000000110;
		15'h2a33: char_row_bitmap <= 16'b0000000000001100;
		15'h2a34: char_row_bitmap <= 16'b0000000000011100;
		15'h2a35: char_row_bitmap <= 16'b0000000000111000;
		15'h2a36: char_row_bitmap <= 16'b0000000001110000;
		15'h2a37: char_row_bitmap <= 16'b0000000001100000;
		15'h2a38: char_row_bitmap <= 16'b0000000011100000;
		15'h2a39: char_row_bitmap <= 16'b0000000111000000;
		15'h2a3a: char_row_bitmap <= 16'b0000001111000000;
		15'h2a3b: char_row_bitmap <= 16'b0000011111100000;
		15'h2a3c: char_row_bitmap <= 16'b0000011001100000;
		15'h2a3d: char_row_bitmap <= 16'b0000111001110000;
		15'h2a3e: char_row_bitmap <= 16'b0001110000111000;
		15'h2a3f: char_row_bitmap <= 16'b0011100000011100;
		15'h2a40: char_row_bitmap <= 16'b0111000000001110;
		15'h2a41: char_row_bitmap <= 16'b0110000000000110;
		15'h2a42: char_row_bitmap <= 16'b1110000000000111;
		15'h2a43: char_row_bitmap <= 16'b1100000000000011;
		15'h2a44: char_row_bitmap <= 16'b0000000000000000;
		15'h2a45: char_row_bitmap <= 16'b0000000000000000;
		15'h2a46: char_row_bitmap <= 16'b0000000000000000;
		15'h2a47: char_row_bitmap <= 16'b0000000000000000;
		15'h2a48: char_row_bitmap <= 16'b0000000000000000;
		15'h2a49: char_row_bitmap <= 16'b0000000000000000;
		15'h2a4a: char_row_bitmap <= 16'b0000000000000000;
		15'h2a4b: char_row_bitmap <= 16'b0000000000000000;
		15'h2a4c: char_row_bitmap <= 16'b0000000000000000;
		15'h2a4d: char_row_bitmap <= 16'b0000000000000000;
		15'h2a4e: char_row_bitmap <= 16'b0000000000000000;
		15'h2a4f: char_row_bitmap <= 16'b0000000000000000;
		15'h2a50: char_row_bitmap <= 16'b0000000000000000;
		15'h2a51: char_row_bitmap <= 16'b0000000000000000;
		15'h2a52: char_row_bitmap <= 16'b0000000000000000;
		15'h2a53: char_row_bitmap <= 16'b0000000000000000;
		15'h2a54: char_row_bitmap <= 16'b0000000000000000;
		15'h2a55: char_row_bitmap <= 16'b0000000000000000;
		15'h2a56: char_row_bitmap <= 16'b0000000000000000;
		15'h2a57: char_row_bitmap <= 16'b0000000000000000;
		15'h2a58: char_row_bitmap <= 16'b0000000000000000;
		15'h2a59: char_row_bitmap <= 16'b0000000000000000;
		15'h2a5a: char_row_bitmap <= 16'b0000000000000000;
		15'h2a5b: char_row_bitmap <= 16'b0000000000000000;
		15'h2a5c: char_row_bitmap <= 16'b0000000000000000;
		15'h2a5d: char_row_bitmap <= 16'b0000000000000000;
		15'h2a5e: char_row_bitmap <= 16'b0000000000000000;
		15'h2a5f: char_row_bitmap <= 16'b0000000000000000;
		15'h2a60: char_row_bitmap <= 16'b0000000000000000;
		15'h2a61: char_row_bitmap <= 16'b0000000000000000;
		15'h2a62: char_row_bitmap <= 16'b0000000000000000;
		15'h2a63: char_row_bitmap <= 16'b0000000000000000;
		15'h2a64: char_row_bitmap <= 16'b0000000000000000;
		15'h2a65: char_row_bitmap <= 16'b0000000000000000;
		15'h2a66: char_row_bitmap <= 16'b0000000000000000;
		15'h2a67: char_row_bitmap <= 16'b0000000000000000;
		15'h2a68: char_row_bitmap <= 16'b0000000000000000;
		15'h2a69: char_row_bitmap <= 16'b0000000000000000;
		15'h2a6a: char_row_bitmap <= 16'b0000000000000000;
		15'h2a6b: char_row_bitmap <= 16'b0000000000000000;
		15'h2a6c: char_row_bitmap <= 16'b1100000000000011;
		15'h2a6d: char_row_bitmap <= 16'b1110000000000111;
		15'h2a6e: char_row_bitmap <= 16'b0110000000000110;
		15'h2a6f: char_row_bitmap <= 16'b0011000000001100;
		15'h2a70: char_row_bitmap <= 16'b0011100000011100;
		15'h2a71: char_row_bitmap <= 16'b0001110000111000;
		15'h2a72: char_row_bitmap <= 16'b0000111001110000;
		15'h2a73: char_row_bitmap <= 16'b0000011001100000;
		15'h2a74: char_row_bitmap <= 16'b0000011111100000;
		15'h2a75: char_row_bitmap <= 16'b0000001111000000;
		15'h2a76: char_row_bitmap <= 16'b0000001111000000;
		15'h2a77: char_row_bitmap <= 16'b0000011111100000;
		15'h2a78: char_row_bitmap <= 16'b0000011001100000;
		15'h2a79: char_row_bitmap <= 16'b0000111001110000;
		15'h2a7a: char_row_bitmap <= 16'b0001110000111000;
		15'h2a7b: char_row_bitmap <= 16'b0011100000011100;
		15'h2a7c: char_row_bitmap <= 16'b0111000000001110;
		15'h2a7d: char_row_bitmap <= 16'b0110000000000110;
		15'h2a7e: char_row_bitmap <= 16'b1110000000000111;
		15'h2a7f: char_row_bitmap <= 16'b1100000000000011;
		15'h2a80: char_row_bitmap <= 16'b0000000000000000;
		15'h2a81: char_row_bitmap <= 16'b0000000000000000;
		15'h2a82: char_row_bitmap <= 16'b0000000000000000;
		15'h2a83: char_row_bitmap <= 16'b0000000000000000;
		15'h2a84: char_row_bitmap <= 16'b0000000000111100;
		15'h2a85: char_row_bitmap <= 16'b0000000000111100;
		15'h2a86: char_row_bitmap <= 16'b0000001000111100;
		15'h2a87: char_row_bitmap <= 16'b0000011000111100;
		15'h2a88: char_row_bitmap <= 16'b0000111000111100;
		15'h2a89: char_row_bitmap <= 16'b0001111001111100;
		15'h2a8a: char_row_bitmap <= 16'b0011111111111000;
		15'h2a8b: char_row_bitmap <= 16'b0111111111111000;
		15'h2a8c: char_row_bitmap <= 16'b0111111111110000;
		15'h2a8d: char_row_bitmap <= 16'b0011111111000000;
		15'h2a8e: char_row_bitmap <= 16'b0001111000000000;
		15'h2a8f: char_row_bitmap <= 16'b0000111000000000;
		15'h2a90: char_row_bitmap <= 16'b0000011000000000;
		15'h2a91: char_row_bitmap <= 16'b0000001000000000;
		15'h2a92: char_row_bitmap <= 16'b0000000000000000;
		15'h2a93: char_row_bitmap <= 16'b0000000000000000;
		15'h2a94: char_row_bitmap <= 16'b0000000111000000;
		15'h2a95: char_row_bitmap <= 16'b0000000011100000;
		15'h2a96: char_row_bitmap <= 16'b0000000001100000;
		15'h2a97: char_row_bitmap <= 16'b0000000001110000;
		15'h2a98: char_row_bitmap <= 16'b0000000000111000;
		15'h2a99: char_row_bitmap <= 16'b0000000000011100;
		15'h2a9a: char_row_bitmap <= 16'b0000000000001110;
		15'h2a9b: char_row_bitmap <= 16'b0000000000000110;
		15'h2a9c: char_row_bitmap <= 16'b0000000000000111;
		15'h2a9d: char_row_bitmap <= 16'b0000000000000011;
		15'h2a9e: char_row_bitmap <= 16'b0000000000000001;
		15'h2a9f: char_row_bitmap <= 16'b0000000000000000;
		15'h2aa0: char_row_bitmap <= 16'b0000000000000000;
		15'h2aa1: char_row_bitmap <= 16'b0000000000000000;
		15'h2aa2: char_row_bitmap <= 16'b0000000000000000;
		15'h2aa3: char_row_bitmap <= 16'b0000000000000000;
		15'h2aa4: char_row_bitmap <= 16'b0000000000000000;
		15'h2aa5: char_row_bitmap <= 16'b0000000000000000;
		15'h2aa6: char_row_bitmap <= 16'b0000000000000000;
		15'h2aa7: char_row_bitmap <= 16'b0000000000000000;
		15'h2aa8: char_row_bitmap <= 16'b0000000000000000;
		15'h2aa9: char_row_bitmap <= 16'b0000000000000000;
		15'h2aaa: char_row_bitmap <= 16'b0000000000000000;
		15'h2aab: char_row_bitmap <= 16'b0000000000000000;
		15'h2aac: char_row_bitmap <= 16'b0000000000000000;
		15'h2aad: char_row_bitmap <= 16'b0000000000000000;
		15'h2aae: char_row_bitmap <= 16'b0000000000000000;
		15'h2aaf: char_row_bitmap <= 16'b0000000000000000;
		15'h2ab0: char_row_bitmap <= 16'b0000000000000000;
		15'h2ab1: char_row_bitmap <= 16'b0000000000000001;
		15'h2ab2: char_row_bitmap <= 16'b0000000000000011;
		15'h2ab3: char_row_bitmap <= 16'b0000000000000111;
		15'h2ab4: char_row_bitmap <= 16'b0000000000000110;
		15'h2ab5: char_row_bitmap <= 16'b0000000000001110;
		15'h2ab6: char_row_bitmap <= 16'b0000000000011100;
		15'h2ab7: char_row_bitmap <= 16'b0000000000111000;
		15'h2ab8: char_row_bitmap <= 16'b0000000001110000;
		15'h2ab9: char_row_bitmap <= 16'b0000000001100000;
		15'h2aba: char_row_bitmap <= 16'b0000000011100000;
		15'h2abb: char_row_bitmap <= 16'b0000000111000000;
		15'h2abc: char_row_bitmap <= 16'b0000000111000000;
		15'h2abd: char_row_bitmap <= 16'b0000000011100000;
		15'h2abe: char_row_bitmap <= 16'b0000000001100000;
		15'h2abf: char_row_bitmap <= 16'b0000000001110000;
		15'h2ac0: char_row_bitmap <= 16'b0000000000111000;
		15'h2ac1: char_row_bitmap <= 16'b0000000000011100;
		15'h2ac2: char_row_bitmap <= 16'b0000000000001110;
		15'h2ac3: char_row_bitmap <= 16'b0000000000000110;
		15'h2ac4: char_row_bitmap <= 16'b0000000000000111;
		15'h2ac5: char_row_bitmap <= 16'b0000000000000011;
		15'h2ac6: char_row_bitmap <= 16'b0000000000000011;
		15'h2ac7: char_row_bitmap <= 16'b0000000000000111;
		15'h2ac8: char_row_bitmap <= 16'b0000000000000110;
		15'h2ac9: char_row_bitmap <= 16'b0000000000001110;
		15'h2aca: char_row_bitmap <= 16'b0000000000011100;
		15'h2acb: char_row_bitmap <= 16'b0000000000111000;
		15'h2acc: char_row_bitmap <= 16'b0000000001110000;
		15'h2acd: char_row_bitmap <= 16'b0000000001100000;
		15'h2ace: char_row_bitmap <= 16'b0000000011100000;
		15'h2acf: char_row_bitmap <= 16'b0000000111000000;
		15'h2ad0: char_row_bitmap <= 16'b0000000000000000;
		15'h2ad1: char_row_bitmap <= 16'b0000000000000000;
		15'h2ad2: char_row_bitmap <= 16'b0000000000000000;
		15'h2ad3: char_row_bitmap <= 16'b0000000000000000;
		15'h2ad4: char_row_bitmap <= 16'b0000000000000000;
		15'h2ad5: char_row_bitmap <= 16'b0000000000000000;
		15'h2ad6: char_row_bitmap <= 16'b0000000000000000;
		15'h2ad7: char_row_bitmap <= 16'b0000000000000000;
		15'h2ad8: char_row_bitmap <= 16'b0000000000000000;
		15'h2ad9: char_row_bitmap <= 16'b1000000000000000;
		15'h2ada: char_row_bitmap <= 16'b1100000000000000;
		15'h2adb: char_row_bitmap <= 16'b1110000000000000;
		15'h2adc: char_row_bitmap <= 16'b0110000000000000;
		15'h2add: char_row_bitmap <= 16'b0111000000000000;
		15'h2ade: char_row_bitmap <= 16'b0011100000000000;
		15'h2adf: char_row_bitmap <= 16'b0001110000000000;
		15'h2ae0: char_row_bitmap <= 16'b0000111000000000;
		15'h2ae1: char_row_bitmap <= 16'b0000011000000000;
		15'h2ae2: char_row_bitmap <= 16'b0000011100000000;
		15'h2ae3: char_row_bitmap <= 16'b0000001110000000;
		15'h2ae4: char_row_bitmap <= 16'b0000000111000000;
		15'h2ae5: char_row_bitmap <= 16'b0000000011100000;
		15'h2ae6: char_row_bitmap <= 16'b0000000001100000;
		15'h2ae7: char_row_bitmap <= 16'b0000000001110000;
		15'h2ae8: char_row_bitmap <= 16'b0000000000111000;
		15'h2ae9: char_row_bitmap <= 16'b0000000000011100;
		15'h2aea: char_row_bitmap <= 16'b0000000000001110;
		15'h2aeb: char_row_bitmap <= 16'b0000000000000110;
		15'h2aec: char_row_bitmap <= 16'b0000000000000111;
		15'h2aed: char_row_bitmap <= 16'b1000000000000011;
		15'h2aee: char_row_bitmap <= 16'b1100000000000001;
		15'h2aef: char_row_bitmap <= 16'b1110000000000000;
		15'h2af0: char_row_bitmap <= 16'b0110000000000000;
		15'h2af1: char_row_bitmap <= 16'b0111000000000000;
		15'h2af2: char_row_bitmap <= 16'b0011100000000000;
		15'h2af3: char_row_bitmap <= 16'b0001110000000000;
		15'h2af4: char_row_bitmap <= 16'b0000111000000000;
		15'h2af5: char_row_bitmap <= 16'b0000011000000000;
		15'h2af6: char_row_bitmap <= 16'b0000011100000000;
		15'h2af7: char_row_bitmap <= 16'b0000001110000000;
		15'h2af8: char_row_bitmap <= 16'b0000000000000000;
		15'h2af9: char_row_bitmap <= 16'b0000000000000000;
		15'h2afa: char_row_bitmap <= 16'b0000000000000000;
		15'h2afb: char_row_bitmap <= 16'b0000000000000000;
		15'h2afc: char_row_bitmap <= 16'b0000000000000000;
		15'h2afd: char_row_bitmap <= 16'b0000000000000000;
		15'h2afe: char_row_bitmap <= 16'b0000000000000000;
		15'h2aff: char_row_bitmap <= 16'b0000000000000000;
		15'h2b00: char_row_bitmap <= 16'b0000000000000000;
		15'h2b01: char_row_bitmap <= 16'b1000000000000001;
		15'h2b02: char_row_bitmap <= 16'b1100000000000011;
		15'h2b03: char_row_bitmap <= 16'b1110000000000111;
		15'h2b04: char_row_bitmap <= 16'b0110000000000110;
		15'h2b05: char_row_bitmap <= 16'b0111000000001110;
		15'h2b06: char_row_bitmap <= 16'b0011100000011100;
		15'h2b07: char_row_bitmap <= 16'b0001110000111000;
		15'h2b08: char_row_bitmap <= 16'b0000111001110000;
		15'h2b09: char_row_bitmap <= 16'b0000011001100000;
		15'h2b0a: char_row_bitmap <= 16'b0000011111100000;
		15'h2b0b: char_row_bitmap <= 16'b0000001111000000;
		15'h2b0c: char_row_bitmap <= 16'b0000000111000000;
		15'h2b0d: char_row_bitmap <= 16'b0000000011100000;
		15'h2b0e: char_row_bitmap <= 16'b0000000001100000;
		15'h2b0f: char_row_bitmap <= 16'b0000000001110000;
		15'h2b10: char_row_bitmap <= 16'b0000000000111000;
		15'h2b11: char_row_bitmap <= 16'b0000000000011100;
		15'h2b12: char_row_bitmap <= 16'b0000000000001110;
		15'h2b13: char_row_bitmap <= 16'b0000000000000110;
		15'h2b14: char_row_bitmap <= 16'b0000000000000111;
		15'h2b15: char_row_bitmap <= 16'b1000000000000011;
		15'h2b16: char_row_bitmap <= 16'b1100000000000011;
		15'h2b17: char_row_bitmap <= 16'b1110000000000111;
		15'h2b18: char_row_bitmap <= 16'b0110000000000110;
		15'h2b19: char_row_bitmap <= 16'b0111000000001110;
		15'h2b1a: char_row_bitmap <= 16'b0011100000011100;
		15'h2b1b: char_row_bitmap <= 16'b0001110000111000;
		15'h2b1c: char_row_bitmap <= 16'b0000111001110000;
		15'h2b1d: char_row_bitmap <= 16'b0000011001100000;
		15'h2b1e: char_row_bitmap <= 16'b0000011111100000;
		15'h2b1f: char_row_bitmap <= 16'b0000001111000000;
		15'h2b20: char_row_bitmap <= 16'b0000001110000000;
		15'h2b21: char_row_bitmap <= 16'b0000011100000000;
		15'h2b22: char_row_bitmap <= 16'b0000011000000000;
		15'h2b23: char_row_bitmap <= 16'b0000111000000000;
		15'h2b24: char_row_bitmap <= 16'b0001110000000000;
		15'h2b25: char_row_bitmap <= 16'b0011100000000000;
		15'h2b26: char_row_bitmap <= 16'b0111000000000000;
		15'h2b27: char_row_bitmap <= 16'b0110000000000000;
		15'h2b28: char_row_bitmap <= 16'b1110000000000000;
		15'h2b29: char_row_bitmap <= 16'b1100000000000000;
		15'h2b2a: char_row_bitmap <= 16'b1000000000000000;
		15'h2b2b: char_row_bitmap <= 16'b0000000000000000;
		15'h2b2c: char_row_bitmap <= 16'b0000000000000000;
		15'h2b2d: char_row_bitmap <= 16'b0000000000000000;
		15'h2b2e: char_row_bitmap <= 16'b0000000000000000;
		15'h2b2f: char_row_bitmap <= 16'b0000000000000000;
		15'h2b30: char_row_bitmap <= 16'b0000000000000000;
		15'h2b31: char_row_bitmap <= 16'b0000000000000000;
		15'h2b32: char_row_bitmap <= 16'b0000000000000000;
		15'h2b33: char_row_bitmap <= 16'b0000000000000000;
		15'h2b34: char_row_bitmap <= 16'b0000001111000000;
		15'h2b35: char_row_bitmap <= 16'b0000011111100000;
		15'h2b36: char_row_bitmap <= 16'b0000011001100000;
		15'h2b37: char_row_bitmap <= 16'b0000111001110000;
		15'h2b38: char_row_bitmap <= 16'b0001110000111000;
		15'h2b39: char_row_bitmap <= 16'b0011100000011100;
		15'h2b3a: char_row_bitmap <= 16'b0111000000001110;
		15'h2b3b: char_row_bitmap <= 16'b0110000000000110;
		15'h2b3c: char_row_bitmap <= 16'b1110000000000111;
		15'h2b3d: char_row_bitmap <= 16'b1100000000000011;
		15'h2b3e: char_row_bitmap <= 16'b1000000000000001;
		15'h2b3f: char_row_bitmap <= 16'b0000000000000000;
		15'h2b40: char_row_bitmap <= 16'b0000000000000000;
		15'h2b41: char_row_bitmap <= 16'b0000000000000000;
		15'h2b42: char_row_bitmap <= 16'b0000000000000000;
		15'h2b43: char_row_bitmap <= 16'b0000000000000000;
		15'h2b44: char_row_bitmap <= 16'b0000000000000000;
		15'h2b45: char_row_bitmap <= 16'b0000000000000000;
		15'h2b46: char_row_bitmap <= 16'b0000000000000000;
		15'h2b47: char_row_bitmap <= 16'b0000000000000000;
		15'h2b48: char_row_bitmap <= 16'b0000001110000000;
		15'h2b49: char_row_bitmap <= 16'b0000011100000000;
		15'h2b4a: char_row_bitmap <= 16'b0000011000000000;
		15'h2b4b: char_row_bitmap <= 16'b0000111000000000;
		15'h2b4c: char_row_bitmap <= 16'b0001110000000000;
		15'h2b4d: char_row_bitmap <= 16'b0011100000000000;
		15'h2b4e: char_row_bitmap <= 16'b0111000000000000;
		15'h2b4f: char_row_bitmap <= 16'b0110000000000000;
		15'h2b50: char_row_bitmap <= 16'b1110000000000000;
		15'h2b51: char_row_bitmap <= 16'b1100000000000001;
		15'h2b52: char_row_bitmap <= 16'b1000000000000011;
		15'h2b53: char_row_bitmap <= 16'b0000000000000111;
		15'h2b54: char_row_bitmap <= 16'b0000000000000110;
		15'h2b55: char_row_bitmap <= 16'b0000000000001110;
		15'h2b56: char_row_bitmap <= 16'b0000000000011100;
		15'h2b57: char_row_bitmap <= 16'b0000000000111000;
		15'h2b58: char_row_bitmap <= 16'b0000000001110000;
		15'h2b59: char_row_bitmap <= 16'b0000000001100000;
		15'h2b5a: char_row_bitmap <= 16'b0000000011100000;
		15'h2b5b: char_row_bitmap <= 16'b0000000111000000;
		15'h2b5c: char_row_bitmap <= 16'b0000001111000000;
		15'h2b5d: char_row_bitmap <= 16'b0000011111100000;
		15'h2b5e: char_row_bitmap <= 16'b0000011001100000;
		15'h2b5f: char_row_bitmap <= 16'b0000111001110000;
		15'h2b60: char_row_bitmap <= 16'b0001110000111000;
		15'h2b61: char_row_bitmap <= 16'b0011100000011100;
		15'h2b62: char_row_bitmap <= 16'b0111000000001110;
		15'h2b63: char_row_bitmap <= 16'b0110000000000110;
		15'h2b64: char_row_bitmap <= 16'b1110000000000111;
		15'h2b65: char_row_bitmap <= 16'b1100000000000011;
		15'h2b66: char_row_bitmap <= 16'b1000000000000011;
		15'h2b67: char_row_bitmap <= 16'b0000000000000111;
		15'h2b68: char_row_bitmap <= 16'b0000000000000110;
		15'h2b69: char_row_bitmap <= 16'b0000000000001110;
		15'h2b6a: char_row_bitmap <= 16'b0000000000011100;
		15'h2b6b: char_row_bitmap <= 16'b0000000000111000;
		15'h2b6c: char_row_bitmap <= 16'b0000000001110000;
		15'h2b6d: char_row_bitmap <= 16'b0000000001100000;
		15'h2b6e: char_row_bitmap <= 16'b0000000011100000;
		15'h2b6f: char_row_bitmap <= 16'b0000000111000000;
		15'h2b70: char_row_bitmap <= 16'b0000001110000000;
		15'h2b71: char_row_bitmap <= 16'b0000011100000000;
		15'h2b72: char_row_bitmap <= 16'b0000011000000000;
		15'h2b73: char_row_bitmap <= 16'b0000111000000000;
		15'h2b74: char_row_bitmap <= 16'b0001110000000000;
		15'h2b75: char_row_bitmap <= 16'b0011100000000000;
		15'h2b76: char_row_bitmap <= 16'b0111000000000000;
		15'h2b77: char_row_bitmap <= 16'b0110000000000000;
		15'h2b78: char_row_bitmap <= 16'b1110000000000000;
		15'h2b79: char_row_bitmap <= 16'b1100000000000000;
		15'h2b7a: char_row_bitmap <= 16'b1100000000000000;
		15'h2b7b: char_row_bitmap <= 16'b1110000000000000;
		15'h2b7c: char_row_bitmap <= 16'b0110000000000000;
		15'h2b7d: char_row_bitmap <= 16'b0111000000000000;
		15'h2b7e: char_row_bitmap <= 16'b0011100000000000;
		15'h2b7f: char_row_bitmap <= 16'b0001110000000000;
		15'h2b80: char_row_bitmap <= 16'b0000111000000000;
		15'h2b81: char_row_bitmap <= 16'b0000011000000000;
		15'h2b82: char_row_bitmap <= 16'b0000011100000000;
		15'h2b83: char_row_bitmap <= 16'b0000001110000000;
		15'h2b84: char_row_bitmap <= 16'b0000001111000000;
		15'h2b85: char_row_bitmap <= 16'b0000011111100000;
		15'h2b86: char_row_bitmap <= 16'b0000011001100000;
		15'h2b87: char_row_bitmap <= 16'b0000111001110000;
		15'h2b88: char_row_bitmap <= 16'b0001110000111000;
		15'h2b89: char_row_bitmap <= 16'b0011100000011100;
		15'h2b8a: char_row_bitmap <= 16'b0111000000001110;
		15'h2b8b: char_row_bitmap <= 16'b0110000000000110;
		15'h2b8c: char_row_bitmap <= 16'b1110000000000111;
		15'h2b8d: char_row_bitmap <= 16'b1100000000000011;
		15'h2b8e: char_row_bitmap <= 16'b1100000000000001;
		15'h2b8f: char_row_bitmap <= 16'b1110000000000000;
		15'h2b90: char_row_bitmap <= 16'b0110000000000000;
		15'h2b91: char_row_bitmap <= 16'b0111000000000000;
		15'h2b92: char_row_bitmap <= 16'b0011100000000000;
		15'h2b93: char_row_bitmap <= 16'b0001110000000000;
		15'h2b94: char_row_bitmap <= 16'b0000111000000000;
		15'h2b95: char_row_bitmap <= 16'b0000011000000000;
		15'h2b96: char_row_bitmap <= 16'b0000011100000000;
		15'h2b97: char_row_bitmap <= 16'b0000001110000000;
		15'h2b98: char_row_bitmap <= 16'b0000001110000000;
		15'h2b99: char_row_bitmap <= 16'b0000011100000000;
		15'h2b9a: char_row_bitmap <= 16'b0000011000000000;
		15'h2b9b: char_row_bitmap <= 16'b0000111000000000;
		15'h2b9c: char_row_bitmap <= 16'b0001110000000000;
		15'h2b9d: char_row_bitmap <= 16'b0011100000000000;
		15'h2b9e: char_row_bitmap <= 16'b0111000000000000;
		15'h2b9f: char_row_bitmap <= 16'b0110000000000000;
		15'h2ba0: char_row_bitmap <= 16'b1110000000000000;
		15'h2ba1: char_row_bitmap <= 16'b1100000000000001;
		15'h2ba2: char_row_bitmap <= 16'b1100000000000011;
		15'h2ba3: char_row_bitmap <= 16'b1110000000000111;
		15'h2ba4: char_row_bitmap <= 16'b0110000000000110;
		15'h2ba5: char_row_bitmap <= 16'b0111000000001110;
		15'h2ba6: char_row_bitmap <= 16'b0011100000011100;
		15'h2ba7: char_row_bitmap <= 16'b0001110000111000;
		15'h2ba8: char_row_bitmap <= 16'b0000111001110000;
		15'h2ba9: char_row_bitmap <= 16'b0000011001100000;
		15'h2baa: char_row_bitmap <= 16'b0000011111100000;
		15'h2bab: char_row_bitmap <= 16'b0000001111000000;
		15'h2bac: char_row_bitmap <= 16'b0000001111000000;
		15'h2bad: char_row_bitmap <= 16'b0000011111100000;
		15'h2bae: char_row_bitmap <= 16'b0000011001100000;
		15'h2baf: char_row_bitmap <= 16'b0000111001110000;
		15'h2bb0: char_row_bitmap <= 16'b0001110000111000;
		15'h2bb1: char_row_bitmap <= 16'b0011100000011100;
		15'h2bb2: char_row_bitmap <= 16'b0111000000001110;
		15'h2bb3: char_row_bitmap <= 16'b0110000000000110;
		15'h2bb4: char_row_bitmap <= 16'b1110000000000111;
		15'h2bb5: char_row_bitmap <= 16'b1100000000000011;
		15'h2bb6: char_row_bitmap <= 16'b1100000000000011;
		15'h2bb7: char_row_bitmap <= 16'b1110000000000111;
		15'h2bb8: char_row_bitmap <= 16'b0110000000000110;
		15'h2bb9: char_row_bitmap <= 16'b0111000000001110;
		15'h2bba: char_row_bitmap <= 16'b0011100000011100;
		15'h2bbb: char_row_bitmap <= 16'b0001110000111000;
		15'h2bbc: char_row_bitmap <= 16'b0000111001110000;
		15'h2bbd: char_row_bitmap <= 16'b0000011001100000;
		15'h2bbe: char_row_bitmap <= 16'b0000011111100000;
		15'h2bbf: char_row_bitmap <= 16'b0000001111000000;
		15'h2bc0: char_row_bitmap <= 16'b0000000110000000;
		15'h2bc1: char_row_bitmap <= 16'b0000000110000000;
		15'h2bc2: char_row_bitmap <= 16'b0001111111111000;
		15'h2bc3: char_row_bitmap <= 16'b0011111111111100;
		15'h2bc4: char_row_bitmap <= 16'b0111111111111110;
		15'h2bc5: char_row_bitmap <= 16'b0111111111111110;
		15'h2bc6: char_row_bitmap <= 16'b0001100110011000;
		15'h2bc7: char_row_bitmap <= 16'b0001100110011000;
		15'h2bc8: char_row_bitmap <= 16'b0001100110011000;
		15'h2bc9: char_row_bitmap <= 16'b0001100110011000;
		15'h2bca: char_row_bitmap <= 16'b0001100110011000;
		15'h2bcb: char_row_bitmap <= 16'b0001100110011000;
		15'h2bcc: char_row_bitmap <= 16'b0001100110011000;
		15'h2bcd: char_row_bitmap <= 16'b0001100110011000;
		15'h2bce: char_row_bitmap <= 16'b0001100000011000;
		15'h2bcf: char_row_bitmap <= 16'b0001100000011000;
		15'h2bd0: char_row_bitmap <= 16'b0001111111111000;
		15'h2bd1: char_row_bitmap <= 16'b0001111111111000;
		15'h2bd2: char_row_bitmap <= 16'b0000000000000000;
		15'h2bd3: char_row_bitmap <= 16'b0000000000000000;
		15'h2bd4: char_row_bitmap <= 16'b0000000110000000;
		15'h2bd5: char_row_bitmap <= 16'b0000000110000000;
		15'h2bd6: char_row_bitmap <= 16'b0001111111111000;
		15'h2bd7: char_row_bitmap <= 16'b0011111111111100;
		15'h2bd8: char_row_bitmap <= 16'b0111111111111110;
		15'h2bd9: char_row_bitmap <= 16'b0111111111111110;
		15'h2bda: char_row_bitmap <= 16'b0001100110011000;
		15'h2bdb: char_row_bitmap <= 16'b0011100110011100;
		15'h2bdc: char_row_bitmap <= 16'b0111000110001110;
		15'h2bdd: char_row_bitmap <= 16'b0110000110000110;
		15'h2bde: char_row_bitmap <= 16'b0110000110000110;
		15'h2bdf: char_row_bitmap <= 16'b0110000110000110;
		15'h2be0: char_row_bitmap <= 16'b0110000110000110;
		15'h2be1: char_row_bitmap <= 16'b0111000110001110;
		15'h2be2: char_row_bitmap <= 16'b0011100000011100;
		15'h2be3: char_row_bitmap <= 16'b0001100000011000;
		15'h2be4: char_row_bitmap <= 16'b0001111111111000;
		15'h2be5: char_row_bitmap <= 16'b0001111111111000;
		15'h2be6: char_row_bitmap <= 16'b0000000000000000;
		15'h2be7: char_row_bitmap <= 16'b0000000000000000;
		15'h2be8: char_row_bitmap <= 16'b0000000000000000;
		15'h2be9: char_row_bitmap <= 16'b0000000000000000;
		15'h2bea: char_row_bitmap <= 16'b0000001111000000;
		15'h2beb: char_row_bitmap <= 16'b0000011111100000;
		15'h2bec: char_row_bitmap <= 16'b0000011111100000;
		15'h2bed: char_row_bitmap <= 16'b0000001111000000;
		15'h2bee: char_row_bitmap <= 16'b0110000110000110;
		15'h2bef: char_row_bitmap <= 16'b0111000110001110;
		15'h2bf0: char_row_bitmap <= 16'b0011111111111100;
		15'h2bf1: char_row_bitmap <= 16'b0001111111111000;
		15'h2bf2: char_row_bitmap <= 16'b0000000110000000;
		15'h2bf3: char_row_bitmap <= 16'b0000001111000000;
		15'h2bf4: char_row_bitmap <= 16'b0000011111100000;
		15'h2bf5: char_row_bitmap <= 16'b0000011001100000;
		15'h2bf6: char_row_bitmap <= 16'b0000011001100000;
		15'h2bf7: char_row_bitmap <= 16'b0000011001100000;
		15'h2bf8: char_row_bitmap <= 16'b0000011001100000;
		15'h2bf9: char_row_bitmap <= 16'b0000011001100000;
		15'h2bfa: char_row_bitmap <= 16'b0000000000000000;
		15'h2bfb: char_row_bitmap <= 16'b0000000000000000;
		15'h2bfc: char_row_bitmap <= 16'b0000000000000000;
		15'h2bfd: char_row_bitmap <= 16'b0000000000000000;
		15'h2bfe: char_row_bitmap <= 16'b0000001111000000;
		15'h2bff: char_row_bitmap <= 16'b0000011111100000;
		15'h2c00: char_row_bitmap <= 16'b0000011111100000;
		15'h2c01: char_row_bitmap <= 16'b0000001111000000;
		15'h2c02: char_row_bitmap <= 16'b0000000110000000;
		15'h2c03: char_row_bitmap <= 16'b0000000110000000;
		15'h2c04: char_row_bitmap <= 16'b0111111111111110;
		15'h2c05: char_row_bitmap <= 16'b0111111111111110;
		15'h2c06: char_row_bitmap <= 16'b0000000110000000;
		15'h2c07: char_row_bitmap <= 16'b0000001111000000;
		15'h2c08: char_row_bitmap <= 16'b0000011111100000;
		15'h2c09: char_row_bitmap <= 16'b0000111001110000;
		15'h2c0a: char_row_bitmap <= 16'b0001110000111000;
		15'h2c0b: char_row_bitmap <= 16'b0011100000011100;
		15'h2c0c: char_row_bitmap <= 16'b0111000000001110;
		15'h2c0d: char_row_bitmap <= 16'b0110000000000110;
		15'h2c0e: char_row_bitmap <= 16'b0000000000000000;
		15'h2c0f: char_row_bitmap <= 16'b0000000000000000;
		15'h2c10: char_row_bitmap <= 16'b0000000000000000;
		15'h2c11: char_row_bitmap <= 16'b0000000000000000;
		15'h2c12: char_row_bitmap <= 16'b0000001111000000;
		15'h2c13: char_row_bitmap <= 16'b0000011111100000;
		15'h2c14: char_row_bitmap <= 16'b0000011111100000;
		15'h2c15: char_row_bitmap <= 16'b0000001111000000;
		15'h2c16: char_row_bitmap <= 16'b0000000110000110;
		15'h2c17: char_row_bitmap <= 16'b0000000110001110;
		15'h2c18: char_row_bitmap <= 16'b0001111111111100;
		15'h2c19: char_row_bitmap <= 16'b0011111111111000;
		15'h2c1a: char_row_bitmap <= 16'b0111000110000000;
		15'h2c1b: char_row_bitmap <= 16'b0110001111000000;
		15'h2c1c: char_row_bitmap <= 16'b0000011111100000;
		15'h2c1d: char_row_bitmap <= 16'b0000011001110000;
		15'h2c1e: char_row_bitmap <= 16'b0000011000111000;
		15'h2c1f: char_row_bitmap <= 16'b0000011000011100;
		15'h2c20: char_row_bitmap <= 16'b0000011000001110;
		15'h2c21: char_row_bitmap <= 16'b0000011000000110;
		15'h2c22: char_row_bitmap <= 16'b0000000000000000;
		15'h2c23: char_row_bitmap <= 16'b0000000000000000;
		15'h2c24: char_row_bitmap <= 16'b0000000000000000;
		15'h2c25: char_row_bitmap <= 16'b0000000000000000;
		15'h2c26: char_row_bitmap <= 16'b0000001111000000;
		15'h2c27: char_row_bitmap <= 16'b0000011111100000;
		15'h2c28: char_row_bitmap <= 16'b0000011111100000;
		15'h2c29: char_row_bitmap <= 16'b0000001111000000;
		15'h2c2a: char_row_bitmap <= 16'b0110000110000000;
		15'h2c2b: char_row_bitmap <= 16'b0111000110000000;
		15'h2c2c: char_row_bitmap <= 16'b0011111111111000;
		15'h2c2d: char_row_bitmap <= 16'b0001111111111100;
		15'h2c2e: char_row_bitmap <= 16'b0000000110001110;
		15'h2c2f: char_row_bitmap <= 16'b0000001111000110;
		15'h2c30: char_row_bitmap <= 16'b0000011111100000;
		15'h2c31: char_row_bitmap <= 16'b0000111001100000;
		15'h2c32: char_row_bitmap <= 16'b0001110001100000;
		15'h2c33: char_row_bitmap <= 16'b0011100001100000;
		15'h2c34: char_row_bitmap <= 16'b0111000001100000;
		15'h2c35: char_row_bitmap <= 16'b0110000001100000;
		15'h2c36: char_row_bitmap <= 16'b0000000000000000;
		15'h2c37: char_row_bitmap <= 16'b0000000000000000;
		15'h2c38: char_row_bitmap <= 16'b0000000000000000;
		15'h2c39: char_row_bitmap <= 16'b0000000000000000;
		15'h2c3a: char_row_bitmap <= 16'b0000000000000000;
		15'h2c3b: char_row_bitmap <= 16'b0000000110000000;
		15'h2c3c: char_row_bitmap <= 16'b0000001111000000;
		15'h2c3d: char_row_bitmap <= 16'b0000011111100000;
		15'h2c3e: char_row_bitmap <= 16'b0000011111100000;
		15'h2c3f: char_row_bitmap <= 16'b0000011111100000;
		15'h2c40: char_row_bitmap <= 16'b0001101111011000;
		15'h2c41: char_row_bitmap <= 16'b0011111111111100;
		15'h2c42: char_row_bitmap <= 16'b0111111111111110;
		15'h2c43: char_row_bitmap <= 16'b0111111111111110;
		15'h2c44: char_row_bitmap <= 16'b0111111111111110;
		15'h2c45: char_row_bitmap <= 16'b0011110110111100;
		15'h2c46: char_row_bitmap <= 16'b0001100110011000;
		15'h2c47: char_row_bitmap <= 16'b0000000110000000;
		15'h2c48: char_row_bitmap <= 16'b0000001111000000;
		15'h2c49: char_row_bitmap <= 16'b0000000000000000;
		15'h2c4a: char_row_bitmap <= 16'b0000000000000000;
		15'h2c4b: char_row_bitmap <= 16'b0000000000000000;
		15'h2c4c: char_row_bitmap <= 16'b0000000000000000;
		15'h2c4d: char_row_bitmap <= 16'b0000000110000000;
		15'h2c4e: char_row_bitmap <= 16'b0000000110000000;
		15'h2c4f: char_row_bitmap <= 16'b0000001111000000;
		15'h2c50: char_row_bitmap <= 16'b0000001111000000;
		15'h2c51: char_row_bitmap <= 16'b0000011111100000;
		15'h2c52: char_row_bitmap <= 16'b0000011111100000;
		15'h2c53: char_row_bitmap <= 16'b0000111111110000;
		15'h2c54: char_row_bitmap <= 16'b0011111111111100;
		15'h2c55: char_row_bitmap <= 16'b0111111111111110;
		15'h2c56: char_row_bitmap <= 16'b0011111111111100;
		15'h2c57: char_row_bitmap <= 16'b0000111111110000;
		15'h2c58: char_row_bitmap <= 16'b0000011111100000;
		15'h2c59: char_row_bitmap <= 16'b0000011111100000;
		15'h2c5a: char_row_bitmap <= 16'b0000001111000000;
		15'h2c5b: char_row_bitmap <= 16'b0000001111000000;
		15'h2c5c: char_row_bitmap <= 16'b0000000110000000;
		15'h2c5d: char_row_bitmap <= 16'b0000000110000000;
		15'h2c5e: char_row_bitmap <= 16'b0000000000000000;
		15'h2c5f: char_row_bitmap <= 16'b0000000000000000;
		15'h2c60: char_row_bitmap <= 16'b0000000000000000;
		15'h2c61: char_row_bitmap <= 16'b0000000000000000;
		15'h2c62: char_row_bitmap <= 16'b0000000000000000;
		15'h2c63: char_row_bitmap <= 16'b0000000000000000;
		15'h2c64: char_row_bitmap <= 16'b0001100000011000;
		15'h2c65: char_row_bitmap <= 16'b0011110000111100;
		15'h2c66: char_row_bitmap <= 16'b0111111001111110;
		15'h2c67: char_row_bitmap <= 16'b0111111111111110;
		15'h2c68: char_row_bitmap <= 16'b0111111111111110;
		15'h2c69: char_row_bitmap <= 16'b0111111111111110;
		15'h2c6a: char_row_bitmap <= 16'b0011111111111100;
		15'h2c6b: char_row_bitmap <= 16'b0001111111111000;
		15'h2c6c: char_row_bitmap <= 16'b0000111111110000;
		15'h2c6d: char_row_bitmap <= 16'b0000011111100000;
		15'h2c6e: char_row_bitmap <= 16'b0000001111000000;
		15'h2c6f: char_row_bitmap <= 16'b0000001111000000;
		15'h2c70: char_row_bitmap <= 16'b0000000110000000;
		15'h2c71: char_row_bitmap <= 16'b0000000000000000;
		15'h2c72: char_row_bitmap <= 16'b0000000000000000;
		15'h2c73: char_row_bitmap <= 16'b0000000000000000;
		15'h2c74: char_row_bitmap <= 16'b0000000000000000;
		15'h2c75: char_row_bitmap <= 16'b0000000000000000;
		15'h2c76: char_row_bitmap <= 16'b0000000110000000;
		15'h2c77: char_row_bitmap <= 16'b0000000110000000;
		15'h2c78: char_row_bitmap <= 16'b0000001111000000;
		15'h2c79: char_row_bitmap <= 16'b0000011111100000;
		15'h2c7a: char_row_bitmap <= 16'b0000011111100000;
		15'h2c7b: char_row_bitmap <= 16'b0000111111110000;
		15'h2c7c: char_row_bitmap <= 16'b0001111111111000;
		15'h2c7d: char_row_bitmap <= 16'b0011111111111100;
		15'h2c7e: char_row_bitmap <= 16'b0111111111111110;
		15'h2c7f: char_row_bitmap <= 16'b0111111111111110;
		15'h2c80: char_row_bitmap <= 16'b0111111111111110;
		15'h2c81: char_row_bitmap <= 16'b0011110110111100;
		15'h2c82: char_row_bitmap <= 16'b0001100110011000;
		15'h2c83: char_row_bitmap <= 16'b0000000110000000;
		15'h2c84: char_row_bitmap <= 16'b0000001111000000;
		15'h2c85: char_row_bitmap <= 16'b0000000000000000;
		15'h2c86: char_row_bitmap <= 16'b0000000000000000;
		15'h2c87: char_row_bitmap <= 16'b0000000000000000;
		15'h2c88: char_row_bitmap <= 16'b0000000000000000;
		15'h2c89: char_row_bitmap <= 16'b0000000000000000;
		15'h2c8a: char_row_bitmap <= 16'b0000000000000000;
		15'h2c8b: char_row_bitmap <= 16'b0000000000000000;
		15'h2c8c: char_row_bitmap <= 16'b0000000000000000;
		15'h2c8d: char_row_bitmap <= 16'b0000000000000000;
		15'h2c8e: char_row_bitmap <= 16'b0000001111000000;
		15'h2c8f: char_row_bitmap <= 16'b0000011111100000;
		15'h2c90: char_row_bitmap <= 16'b0000111001110000;
		15'h2c91: char_row_bitmap <= 16'b0000110000110000;
		15'h2c92: char_row_bitmap <= 16'b0000110000110000;
		15'h2c93: char_row_bitmap <= 16'b0000111001110000;
		15'h2c94: char_row_bitmap <= 16'b0000011111100000;
		15'h2c95: char_row_bitmap <= 16'b0000001111000000;
		15'h2c96: char_row_bitmap <= 16'b0000000000000000;
		15'h2c97: char_row_bitmap <= 16'b0000000000000000;
		15'h2c98: char_row_bitmap <= 16'b0000000000000000;
		15'h2c99: char_row_bitmap <= 16'b0000000000000000;
		15'h2c9a: char_row_bitmap <= 16'b0000000000000000;
		15'h2c9b: char_row_bitmap <= 16'b0000000000000000;
		15'h2c9c: char_row_bitmap <= 16'b0000000000000000;
		15'h2c9d: char_row_bitmap <= 16'b0000000000000000;
		15'h2c9e: char_row_bitmap <= 16'b0000000000000000;
		15'h2c9f: char_row_bitmap <= 16'b0000000000000000;
		15'h2ca0: char_row_bitmap <= 16'b0000000000000000;
		15'h2ca1: char_row_bitmap <= 16'b0000000000000000;
		15'h2ca2: char_row_bitmap <= 16'b0000001111000000;
		15'h2ca3: char_row_bitmap <= 16'b0000011111100000;
		15'h2ca4: char_row_bitmap <= 16'b0000111111110000;
		15'h2ca5: char_row_bitmap <= 16'b0000111111110000;
		15'h2ca6: char_row_bitmap <= 16'b0000111111110000;
		15'h2ca7: char_row_bitmap <= 16'b0000111111110000;
		15'h2ca8: char_row_bitmap <= 16'b0000011111100000;
		15'h2ca9: char_row_bitmap <= 16'b0000001111000000;
		15'h2caa: char_row_bitmap <= 16'b0000000000000000;
		15'h2cab: char_row_bitmap <= 16'b0000000000000000;
		15'h2cac: char_row_bitmap <= 16'b0000000000000000;
		15'h2cad: char_row_bitmap <= 16'b0000000000000000;
		15'h2cae: char_row_bitmap <= 16'b0000000000000000;
		15'h2caf: char_row_bitmap <= 16'b0000000000000000;
		15'h2cb0: char_row_bitmap <= 16'b0000000000000000;
		15'h2cb1: char_row_bitmap <= 16'b0000000000000000;
		15'h2cb2: char_row_bitmap <= 16'b0000000000000000;
		15'h2cb3: char_row_bitmap <= 16'b0000000000000000;
		15'h2cb4: char_row_bitmap <= 16'b0000011111100000;
		15'h2cb5: char_row_bitmap <= 16'b0001111111111000;
		15'h2cb6: char_row_bitmap <= 16'b0001110000111000;
		15'h2cb7: char_row_bitmap <= 16'b0011100000011100;
		15'h2cb8: char_row_bitmap <= 16'b0011000000001100;
		15'h2cb9: char_row_bitmap <= 16'b0011000000001100;
		15'h2cba: char_row_bitmap <= 16'b0011000000001100;
		15'h2cbb: char_row_bitmap <= 16'b0011000000001100;
		15'h2cbc: char_row_bitmap <= 16'b0011100000011100;
		15'h2cbd: char_row_bitmap <= 16'b0001110000111000;
		15'h2cbe: char_row_bitmap <= 16'b0001111111111000;
		15'h2cbf: char_row_bitmap <= 16'b0000011111100000;
		15'h2cc0: char_row_bitmap <= 16'b0000000000000000;
		15'h2cc1: char_row_bitmap <= 16'b0000000000000000;
		15'h2cc2: char_row_bitmap <= 16'b0000000000000000;
		15'h2cc3: char_row_bitmap <= 16'b0000000000000000;
		15'h2cc4: char_row_bitmap <= 16'b0000000000000000;
		15'h2cc5: char_row_bitmap <= 16'b0000000000000000;
		15'h2cc6: char_row_bitmap <= 16'b0000000000000000;
		15'h2cc7: char_row_bitmap <= 16'b0000000000000000;
		15'h2cc8: char_row_bitmap <= 16'b0000011111100000;
		15'h2cc9: char_row_bitmap <= 16'b0001111111111000;
		15'h2cca: char_row_bitmap <= 16'b0001111111111000;
		15'h2ccb: char_row_bitmap <= 16'b0011111111111100;
		15'h2ccc: char_row_bitmap <= 16'b0011111111111100;
		15'h2ccd: char_row_bitmap <= 16'b0011111111111100;
		15'h2cce: char_row_bitmap <= 16'b0011111111111100;
		15'h2ccf: char_row_bitmap <= 16'b0011111111111100;
		15'h2cd0: char_row_bitmap <= 16'b0011111111111100;
		15'h2cd1: char_row_bitmap <= 16'b0001111111111000;
		15'h2cd2: char_row_bitmap <= 16'b0001111111111000;
		15'h2cd3: char_row_bitmap <= 16'b0000011111100000;
		15'h2cd4: char_row_bitmap <= 16'b0000000000000000;
		15'h2cd5: char_row_bitmap <= 16'b0000000000000000;
		15'h2cd6: char_row_bitmap <= 16'b0000000000000000;
		15'h2cd7: char_row_bitmap <= 16'b0000000000000000;
		15'h2cd8: char_row_bitmap <= 16'b0000000000000000;
		15'h2cd9: char_row_bitmap <= 16'b0000000000000000;
		15'h2cda: char_row_bitmap <= 16'b0000000000000000;
		15'h2cdb: char_row_bitmap <= 16'b0000000100000000;
		15'h2cdc: char_row_bitmap <= 16'b0000000100000000;
		15'h2cdd: char_row_bitmap <= 16'b0000001110000000;
		15'h2cde: char_row_bitmap <= 16'b0000001110000000;
		15'h2cdf: char_row_bitmap <= 16'b0000001110000000;
		15'h2ce0: char_row_bitmap <= 16'b0111111111111100;
		15'h2ce1: char_row_bitmap <= 16'b0011111111111000;
		15'h2ce2: char_row_bitmap <= 16'b0000111111100000;
		15'h2ce3: char_row_bitmap <= 16'b0000011111000000;
		15'h2ce4: char_row_bitmap <= 16'b0000111111100000;
		15'h2ce5: char_row_bitmap <= 16'b0000111011100000;
		15'h2ce6: char_row_bitmap <= 16'b0001100000110000;
		15'h2ce7: char_row_bitmap <= 16'b0001000000010000;
		15'h2ce8: char_row_bitmap <= 16'b0000000000000000;
		15'h2ce9: char_row_bitmap <= 16'b0000000000000000;
		15'h2cea: char_row_bitmap <= 16'b0000000000000000;
		15'h2ceb: char_row_bitmap <= 16'b0000000000000000;
		15'h2cec: char_row_bitmap <= 16'b0000000000000000;
		15'h2ced: char_row_bitmap <= 16'b0000000000000000;
		15'h2cee: char_row_bitmap <= 16'b0000000000000000;
		15'h2cef: char_row_bitmap <= 16'b0000000000000000;
		15'h2cf0: char_row_bitmap <= 16'b0001110000000000;
		15'h2cf1: char_row_bitmap <= 16'b0000011110000000;
		15'h2cf2: char_row_bitmap <= 16'b0000001111000000;
		15'h2cf3: char_row_bitmap <= 16'b0000000111100000;
		15'h2cf4: char_row_bitmap <= 16'b0000000011110000;
		15'h2cf5: char_row_bitmap <= 16'b0000000011110000;
		15'h2cf6: char_row_bitmap <= 16'b0000000011111000;
		15'h2cf7: char_row_bitmap <= 16'b0000000011111000;
		15'h2cf8: char_row_bitmap <= 16'b0000000011110000;
		15'h2cf9: char_row_bitmap <= 16'b0000000011110000;
		15'h2cfa: char_row_bitmap <= 16'b0000000111100000;
		15'h2cfb: char_row_bitmap <= 16'b0000001111000000;
		15'h2cfc: char_row_bitmap <= 16'b0000011110000000;
		15'h2cfd: char_row_bitmap <= 16'b0001110000000000;
		15'h2cfe: char_row_bitmap <= 16'b0000000000000000;
		15'h2cff: char_row_bitmap <= 16'b0000000000000000;
		15'h2d00: char_row_bitmap <= 16'b0000000000000000;
		15'h2d01: char_row_bitmap <= 16'b0000000000000000;
		15'h2d02: char_row_bitmap <= 16'b0000011111100000;
		15'h2d03: char_row_bitmap <= 16'b0001111111111000;
		15'h2d04: char_row_bitmap <= 16'b0011111111111100;
		15'h2d05: char_row_bitmap <= 16'b0011111111111100;
		15'h2d06: char_row_bitmap <= 16'b0111100110011110;
		15'h2d07: char_row_bitmap <= 16'b0111100110011110;
		15'h2d08: char_row_bitmap <= 16'b0111100110011110;
		15'h2d09: char_row_bitmap <= 16'b0111111111111110;
		15'h2d0a: char_row_bitmap <= 16'b0111111111111110;
		15'h2d0b: char_row_bitmap <= 16'b0111111111111110;
		15'h2d0c: char_row_bitmap <= 16'b0110111111110110;
		15'h2d0d: char_row_bitmap <= 16'b0111001111001110;
		15'h2d0e: char_row_bitmap <= 16'b0011110000111100;
		15'h2d0f: char_row_bitmap <= 16'b0011111111111100;
		15'h2d10: char_row_bitmap <= 16'b0001111111111000;
		15'h2d11: char_row_bitmap <= 16'b0000011111100000;
		15'h2d12: char_row_bitmap <= 16'b0000000000000000;
		15'h2d13: char_row_bitmap <= 16'b0000000000000000;
		15'h2d14: char_row_bitmap <= 16'b0000000000000000;
		15'h2d15: char_row_bitmap <= 16'b0000000000000000;
		15'h2d16: char_row_bitmap <= 16'b0000011111100000;
		15'h2d17: char_row_bitmap <= 16'b0001111111111000;
		15'h2d18: char_row_bitmap <= 16'b0011111111111100;
		15'h2d19: char_row_bitmap <= 16'b0011111111111100;
		15'h2d1a: char_row_bitmap <= 16'b0111100110011110;
		15'h2d1b: char_row_bitmap <= 16'b0111100110011110;
		15'h2d1c: char_row_bitmap <= 16'b0111100110011110;
		15'h2d1d: char_row_bitmap <= 16'b0111111111111110;
		15'h2d1e: char_row_bitmap <= 16'b0111111111111110;
		15'h2d1f: char_row_bitmap <= 16'b0111111111111110;
		15'h2d20: char_row_bitmap <= 16'b0110000000000110;
		15'h2d21: char_row_bitmap <= 16'b0111111111111110;
		15'h2d22: char_row_bitmap <= 16'b0011111111111100;
		15'h2d23: char_row_bitmap <= 16'b0011111111111100;
		15'h2d24: char_row_bitmap <= 16'b0001111111111000;
		15'h2d25: char_row_bitmap <= 16'b0000011111100000;
		15'h2d26: char_row_bitmap <= 16'b0000000000000000;
		15'h2d27: char_row_bitmap <= 16'b0000000000000000;
		15'h2d28: char_row_bitmap <= 16'b0000000000000000;
		15'h2d29: char_row_bitmap <= 16'b0000000000000000;
		15'h2d2a: char_row_bitmap <= 16'b0000011111100000;
		15'h2d2b: char_row_bitmap <= 16'b0001111111111000;
		15'h2d2c: char_row_bitmap <= 16'b0011111111111100;
		15'h2d2d: char_row_bitmap <= 16'b0011111111111100;
		15'h2d2e: char_row_bitmap <= 16'b0111100110011110;
		15'h2d2f: char_row_bitmap <= 16'b0111100110011110;
		15'h2d30: char_row_bitmap <= 16'b0111100110011110;
		15'h2d31: char_row_bitmap <= 16'b0111111111111110;
		15'h2d32: char_row_bitmap <= 16'b0111110000111110;
		15'h2d33: char_row_bitmap <= 16'b0111001111001110;
		15'h2d34: char_row_bitmap <= 16'b0110111111110110;
		15'h2d35: char_row_bitmap <= 16'b0111111111111110;
		15'h2d36: char_row_bitmap <= 16'b0011111111111100;
		15'h2d37: char_row_bitmap <= 16'b0011111111111100;
		15'h2d38: char_row_bitmap <= 16'b0001111111111000;
		15'h2d39: char_row_bitmap <= 16'b0000011111100000;
		15'h2d3a: char_row_bitmap <= 16'b0000000000000000;
		15'h2d3b: char_row_bitmap <= 16'b0000000000000000;
		15'h2d3c: char_row_bitmap <= 16'b0000000000000000;
		15'h2d3d: char_row_bitmap <= 16'b0000000000000000;
		15'h2d3e: char_row_bitmap <= 16'b0000011111100000;
		15'h2d3f: char_row_bitmap <= 16'b0001111111111000;
		15'h2d40: char_row_bitmap <= 16'b0011111111111100;
		15'h2d41: char_row_bitmap <= 16'b0011111111111100;
		15'h2d42: char_row_bitmap <= 16'b0111100111111110;
		15'h2d43: char_row_bitmap <= 16'b0111100110001110;
		15'h2d44: char_row_bitmap <= 16'b0111100111111110;
		15'h2d45: char_row_bitmap <= 16'b0111111111111110;
		15'h2d46: char_row_bitmap <= 16'b0111111111111110;
		15'h2d47: char_row_bitmap <= 16'b0111111111111110;
		15'h2d48: char_row_bitmap <= 16'b0110111111110110;
		15'h2d49: char_row_bitmap <= 16'b0111001111001110;
		15'h2d4a: char_row_bitmap <= 16'b0011110000111100;
		15'h2d4b: char_row_bitmap <= 16'b0011111111111100;
		15'h2d4c: char_row_bitmap <= 16'b0001111111111000;
		15'h2d4d: char_row_bitmap <= 16'b0000011111100000;
		15'h2d4e: char_row_bitmap <= 16'b0000000000000000;
		15'h2d4f: char_row_bitmap <= 16'b0000000000000000;
		15'h2d50: char_row_bitmap <= 16'b0000000000000000;
		15'h2d51: char_row_bitmap <= 16'b0000000000000000;
		15'h2d52: char_row_bitmap <= 16'b0000011111100000;
		15'h2d53: char_row_bitmap <= 16'b0001111111111000;
		15'h2d54: char_row_bitmap <= 16'b0011111111111100;
		15'h2d55: char_row_bitmap <= 16'b0011111111111100;
		15'h2d56: char_row_bitmap <= 16'b0111100110011110;
		15'h2d57: char_row_bitmap <= 16'b0111100110011110;
		15'h2d58: char_row_bitmap <= 16'b0111100110011110;
		15'h2d59: char_row_bitmap <= 16'b0111111111111110;
		15'h2d5a: char_row_bitmap <= 16'b0110111111110110;
		15'h2d5b: char_row_bitmap <= 16'b0111000000001110;
		15'h2d5c: char_row_bitmap <= 16'b0111101011011110;
		15'h2d5d: char_row_bitmap <= 16'b0111101101011110;
		15'h2d5e: char_row_bitmap <= 16'b0011101111011100;
		15'h2d5f: char_row_bitmap <= 16'b0011110000111100;
		15'h2d60: char_row_bitmap <= 16'b0001111111111000;
		15'h2d61: char_row_bitmap <= 16'b0000011111100000;
		15'h2d62: char_row_bitmap <= 16'b0000000000000000;
		15'h2d63: char_row_bitmap <= 16'b0000000000000000;
		15'h2d64: char_row_bitmap <= 16'b0000000000000000;
		15'h2d65: char_row_bitmap <= 16'b0000000000000000;
		15'h2d66: char_row_bitmap <= 16'b0000011111100000;
		15'h2d67: char_row_bitmap <= 16'b0001100000011000;
		15'h2d68: char_row_bitmap <= 16'b0010000000000100;
		15'h2d69: char_row_bitmap <= 16'b0010000000000100;
		15'h2d6a: char_row_bitmap <= 16'b0100011001100010;
		15'h2d6b: char_row_bitmap <= 16'b0100011001100010;
		15'h2d6c: char_row_bitmap <= 16'b0100011001100010;
		15'h2d6d: char_row_bitmap <= 16'b0100000000000010;
		15'h2d6e: char_row_bitmap <= 16'b0100000000000010;
		15'h2d6f: char_row_bitmap <= 16'b0100000000000010;
		15'h2d70: char_row_bitmap <= 16'b0101000000001010;
		15'h2d71: char_row_bitmap <= 16'b0100110000110010;
		15'h2d72: char_row_bitmap <= 16'b0010001111000100;
		15'h2d73: char_row_bitmap <= 16'b0010000000000100;
		15'h2d74: char_row_bitmap <= 16'b0001100000011000;
		15'h2d75: char_row_bitmap <= 16'b0000011111100000;
		15'h2d76: char_row_bitmap <= 16'b0000000000000000;
		15'h2d77: char_row_bitmap <= 16'b0000000000000000;
		15'h2d78: char_row_bitmap <= 16'b0000000000000000;
		15'h2d79: char_row_bitmap <= 16'b0000000000000000;
		15'h2d7a: char_row_bitmap <= 16'b0000011111100000;
		15'h2d7b: char_row_bitmap <= 16'b0001100000011000;
		15'h2d7c: char_row_bitmap <= 16'b0010000000000100;
		15'h2d7d: char_row_bitmap <= 16'b0010000000000100;
		15'h2d7e: char_row_bitmap <= 16'b0100011001100010;
		15'h2d7f: char_row_bitmap <= 16'b0100011001100010;
		15'h2d80: char_row_bitmap <= 16'b0100011001100010;
		15'h2d81: char_row_bitmap <= 16'b0100000000000010;
		15'h2d82: char_row_bitmap <= 16'b0100000000000010;
		15'h2d83: char_row_bitmap <= 16'b0100000000000010;
		15'h2d84: char_row_bitmap <= 16'b0101111111111010;
		15'h2d85: char_row_bitmap <= 16'b0100000000000010;
		15'h2d86: char_row_bitmap <= 16'b0010000000000100;
		15'h2d87: char_row_bitmap <= 16'b0010000000000100;
		15'h2d88: char_row_bitmap <= 16'b0001100000011000;
		15'h2d89: char_row_bitmap <= 16'b0000011111100000;
		15'h2d8a: char_row_bitmap <= 16'b0000000000000000;
		15'h2d8b: char_row_bitmap <= 16'b0000000000000000;
		15'h2d8c: char_row_bitmap <= 16'b0000000000000000;
		15'h2d8d: char_row_bitmap <= 16'b0000000000000000;
		15'h2d8e: char_row_bitmap <= 16'b0000011111100000;
		15'h2d8f: char_row_bitmap <= 16'b0001100000011000;
		15'h2d90: char_row_bitmap <= 16'b0010000000000100;
		15'h2d91: char_row_bitmap <= 16'b0010000000000100;
		15'h2d92: char_row_bitmap <= 16'b0100011001100010;
		15'h2d93: char_row_bitmap <= 16'b0100011001100010;
		15'h2d94: char_row_bitmap <= 16'b0100011001100010;
		15'h2d95: char_row_bitmap <= 16'b0100000000000010;
		15'h2d96: char_row_bitmap <= 16'b0100001111000010;
		15'h2d97: char_row_bitmap <= 16'b0100110000110010;
		15'h2d98: char_row_bitmap <= 16'b0101000000001010;
		15'h2d99: char_row_bitmap <= 16'b0100000000000010;
		15'h2d9a: char_row_bitmap <= 16'b0010000000000100;
		15'h2d9b: char_row_bitmap <= 16'b0010000000000100;
		15'h2d9c: char_row_bitmap <= 16'b0001100000011000;
		15'h2d9d: char_row_bitmap <= 16'b0000011111100000;
		15'h2d9e: char_row_bitmap <= 16'b0000000000000000;
		15'h2d9f: char_row_bitmap <= 16'b0000000000000000;
		15'h2da0: char_row_bitmap <= 16'b0000000000000000;
		15'h2da1: char_row_bitmap <= 16'b0000000000000000;
		15'h2da2: char_row_bitmap <= 16'b0000011111100000;
		15'h2da3: char_row_bitmap <= 16'b0001100000011000;
		15'h2da4: char_row_bitmap <= 16'b0010000000000100;
		15'h2da5: char_row_bitmap <= 16'b0010000000000100;
		15'h2da6: char_row_bitmap <= 16'b0100011000000010;
		15'h2da7: char_row_bitmap <= 16'b0100011001110010;
		15'h2da8: char_row_bitmap <= 16'b0100011000000010;
		15'h2da9: char_row_bitmap <= 16'b0100000000000010;
		15'h2daa: char_row_bitmap <= 16'b0100000000000010;
		15'h2dab: char_row_bitmap <= 16'b0100000000000010;
		15'h2dac: char_row_bitmap <= 16'b0101000000001010;
		15'h2dad: char_row_bitmap <= 16'b0100110000110010;
		15'h2dae: char_row_bitmap <= 16'b0010001111000100;
		15'h2daf: char_row_bitmap <= 16'b0010000000000100;
		15'h2db0: char_row_bitmap <= 16'b0001100000011000;
		15'h2db1: char_row_bitmap <= 16'b0000011111100000;
		15'h2db2: char_row_bitmap <= 16'b0000000000000000;
		15'h2db3: char_row_bitmap <= 16'b0000000000000000;
		15'h2db4: char_row_bitmap <= 16'b0000000000000000;
		15'h2db5: char_row_bitmap <= 16'b0000000000000000;
		15'h2db6: char_row_bitmap <= 16'b0000011111100000;
		15'h2db7: char_row_bitmap <= 16'b0001100000011000;
		15'h2db8: char_row_bitmap <= 16'b0010000000000100;
		15'h2db9: char_row_bitmap <= 16'b0010000000000100;
		15'h2dba: char_row_bitmap <= 16'b0100011001100010;
		15'h2dbb: char_row_bitmap <= 16'b0100011001100010;
		15'h2dbc: char_row_bitmap <= 16'b0100011001100010;
		15'h2dbd: char_row_bitmap <= 16'b0100000000000010;
		15'h2dbe: char_row_bitmap <= 16'b0101000000001010;
		15'h2dbf: char_row_bitmap <= 16'b0100111111110010;
		15'h2dc0: char_row_bitmap <= 16'b0100010100100010;
		15'h2dc1: char_row_bitmap <= 16'b0100010010100010;
		15'h2dc2: char_row_bitmap <= 16'b0010010000100100;
		15'h2dc3: char_row_bitmap <= 16'b0010001111000100;
		15'h2dc4: char_row_bitmap <= 16'b0001100000011000;
		15'h2dc5: char_row_bitmap <= 16'b0000011111100000;
		15'h2dc6: char_row_bitmap <= 16'b0000000000000000;
		15'h2dc7: char_row_bitmap <= 16'b0000000000000000;
		15'h2dc8: char_row_bitmap <= 16'b0000000000000000;
		15'h2dc9: char_row_bitmap <= 16'b0000000000000000;
		15'h2dca: char_row_bitmap <= 16'b0000000110000000;
		15'h2dcb: char_row_bitmap <= 16'b0000001111000000;
		15'h2dcc: char_row_bitmap <= 16'b0000011111100000;
		15'h2dcd: char_row_bitmap <= 16'b0000111111110000;
		15'h2dce: char_row_bitmap <= 16'b0001110110111000;
		15'h2dcf: char_row_bitmap <= 16'b0001100110011000;
		15'h2dd0: char_row_bitmap <= 16'b0000000110000000;
		15'h2dd1: char_row_bitmap <= 16'b0000000110000000;
		15'h2dd2: char_row_bitmap <= 16'b0000000110000000;
		15'h2dd3: char_row_bitmap <= 16'b0000000110000000;
		15'h2dd4: char_row_bitmap <= 16'b0000000110000000;
		15'h2dd5: char_row_bitmap <= 16'b0000000110000000;
		15'h2dd6: char_row_bitmap <= 16'b0000000110000000;
		15'h2dd7: char_row_bitmap <= 16'b0000000110000000;
		15'h2dd8: char_row_bitmap <= 16'b0000000110000000;
		15'h2dd9: char_row_bitmap <= 16'b0000000110000000;
		15'h2dda: char_row_bitmap <= 16'b0000000110000000;
		15'h2ddb: char_row_bitmap <= 16'b0000000110000000;
		15'h2ddc: char_row_bitmap <= 16'b0000000000000000;
		15'h2ddd: char_row_bitmap <= 16'b0000000000000000;
		15'h2dde: char_row_bitmap <= 16'b0000000000000000;
		15'h2ddf: char_row_bitmap <= 16'b0000000000000000;
		15'h2de0: char_row_bitmap <= 16'b0000000000000000;
		15'h2de1: char_row_bitmap <= 16'b0000001100000000;
		15'h2de2: char_row_bitmap <= 16'b0000001110000000;
		15'h2de3: char_row_bitmap <= 16'b0000000111000000;
		15'h2de4: char_row_bitmap <= 16'b0000000011100000;
		15'h2de5: char_row_bitmap <= 16'b1111111111110000;
		15'h2de6: char_row_bitmap <= 16'b1111111111110000;
		15'h2de7: char_row_bitmap <= 16'b0000000011100000;
		15'h2de8: char_row_bitmap <= 16'b0000000111000000;
		15'h2de9: char_row_bitmap <= 16'b0000001110000000;
		15'h2dea: char_row_bitmap <= 16'b0000001100000000;
		15'h2deb: char_row_bitmap <= 16'b0000000000000000;
		15'h2dec: char_row_bitmap <= 16'b0000000000000000;
		15'h2ded: char_row_bitmap <= 16'b0000000000000000;
		15'h2dee: char_row_bitmap <= 16'b0000000000000000;
		15'h2def: char_row_bitmap <= 16'b0000000000000000;
		15'h2df0: char_row_bitmap <= 16'b0000000110000000;
		15'h2df1: char_row_bitmap <= 16'b0000000110000000;
		15'h2df2: char_row_bitmap <= 16'b0000000110000000;
		15'h2df3: char_row_bitmap <= 16'b0000000110000000;
		15'h2df4: char_row_bitmap <= 16'b0000000110000000;
		15'h2df5: char_row_bitmap <= 16'b0000000110000000;
		15'h2df6: char_row_bitmap <= 16'b0000000110000000;
		15'h2df7: char_row_bitmap <= 16'b0000000110000000;
		15'h2df8: char_row_bitmap <= 16'b0000000110000000;
		15'h2df9: char_row_bitmap <= 16'b0000000110000000;
		15'h2dfa: char_row_bitmap <= 16'b0000000110000000;
		15'h2dfb: char_row_bitmap <= 16'b0000000110000000;
		15'h2dfc: char_row_bitmap <= 16'b0001100110011000;
		15'h2dfd: char_row_bitmap <= 16'b0001110110111000;
		15'h2dfe: char_row_bitmap <= 16'b0000111111110000;
		15'h2dff: char_row_bitmap <= 16'b0000011111100000;
		15'h2e00: char_row_bitmap <= 16'b0000001111000000;
		15'h2e01: char_row_bitmap <= 16'b0000000110000000;
		15'h2e02: char_row_bitmap <= 16'b0000000000000000;
		15'h2e03: char_row_bitmap <= 16'b0000000000000000;
		15'h2e04: char_row_bitmap <= 16'b0000000000000000;
		15'h2e05: char_row_bitmap <= 16'b0000000000000000;
		15'h2e06: char_row_bitmap <= 16'b0000000000000000;
		15'h2e07: char_row_bitmap <= 16'b0000000000000000;
		15'h2e08: char_row_bitmap <= 16'b0000000000000000;
		15'h2e09: char_row_bitmap <= 16'b0000001100000000;
		15'h2e0a: char_row_bitmap <= 16'b0000011100000000;
		15'h2e0b: char_row_bitmap <= 16'b0000111000000000;
		15'h2e0c: char_row_bitmap <= 16'b0001110000000000;
		15'h2e0d: char_row_bitmap <= 16'b0011111111111111;
		15'h2e0e: char_row_bitmap <= 16'b0011111111111111;
		15'h2e0f: char_row_bitmap <= 16'b0001110000000000;
		15'h2e10: char_row_bitmap <= 16'b0000111000000000;
		15'h2e11: char_row_bitmap <= 16'b0000011100000000;
		15'h2e12: char_row_bitmap <= 16'b0000001100000000;
		15'h2e13: char_row_bitmap <= 16'b0000000000000000;
		15'h2e14: char_row_bitmap <= 16'b0000000000000000;
		15'h2e15: char_row_bitmap <= 16'b0000000000000000;
		15'h2e16: char_row_bitmap <= 16'b0000000000000000;
		15'h2e17: char_row_bitmap <= 16'b0000000000000000;
		15'h2e18: char_row_bitmap <= 16'b0000000000000000;
		15'h2e19: char_row_bitmap <= 16'b0000000000000000;
		15'h2e1a: char_row_bitmap <= 16'b0000000000000000;
		15'h2e1b: char_row_bitmap <= 16'b0000000000000000;
		15'h2e1c: char_row_bitmap <= 16'b0000000011000000;
		15'h2e1d: char_row_bitmap <= 16'b0000000011000000;
		15'h2e1e: char_row_bitmap <= 16'b0000000111100000;
		15'h2e1f: char_row_bitmap <= 16'b0000000111100000;
		15'h2e20: char_row_bitmap <= 16'b0000001100110000;
		15'h2e21: char_row_bitmap <= 16'b0000001100111000;
		15'h2e22: char_row_bitmap <= 16'b0000011000011111;
		15'h2e23: char_row_bitmap <= 16'b0001111000001111;
		15'h2e24: char_row_bitmap <= 16'b0011110000000000;
		15'h2e25: char_row_bitmap <= 16'b0111000000000000;
		15'h2e26: char_row_bitmap <= 16'b0110000000000000;
		15'h2e27: char_row_bitmap <= 16'b1110000000000000;
		15'h2e28: char_row_bitmap <= 16'b1100000000000000;
		15'h2e29: char_row_bitmap <= 16'b1100000000000000;
		15'h2e2a: char_row_bitmap <= 16'b0000000000000000;
		15'h2e2b: char_row_bitmap <= 16'b0000000000000000;
		15'h2e2c: char_row_bitmap <= 16'b0000000000000000;
		15'h2e2d: char_row_bitmap <= 16'b0000000000000000;
		15'h2e2e: char_row_bitmap <= 16'b1100000000000000;
		15'h2e2f: char_row_bitmap <= 16'b1100000000000000;
		15'h2e30: char_row_bitmap <= 16'b1110000000000000;
		15'h2e31: char_row_bitmap <= 16'b0110000000000000;
		15'h2e32: char_row_bitmap <= 16'b0111000000000000;
		15'h2e33: char_row_bitmap <= 16'b0011110000000000;
		15'h2e34: char_row_bitmap <= 16'b0001111000001111;
		15'h2e35: char_row_bitmap <= 16'b0000011000011111;
		15'h2e36: char_row_bitmap <= 16'b0000001100111000;
		15'h2e37: char_row_bitmap <= 16'b0000001100110000;
		15'h2e38: char_row_bitmap <= 16'b0000000111100000;
		15'h2e39: char_row_bitmap <= 16'b0000000111100000;
		15'h2e3a: char_row_bitmap <= 16'b0000000011000000;
		15'h2e3b: char_row_bitmap <= 16'b0000000011000000;
		15'h2e3c: char_row_bitmap <= 16'b0000000000000000;
		15'h2e3d: char_row_bitmap <= 16'b0000000000000000;
		15'h2e3e: char_row_bitmap <= 16'b0000000000000000;
		15'h2e3f: char_row_bitmap <= 16'b0000000000000000;
		15'h2e40: char_row_bitmap <= 16'b0000000000000000;
		15'h2e41: char_row_bitmap <= 16'b0000000000000000;
		15'h2e42: char_row_bitmap <= 16'b0000000000000000;
		15'h2e43: char_row_bitmap <= 16'b0000000000000000;
		15'h2e44: char_row_bitmap <= 16'b0000000000000000;
		15'h2e45: char_row_bitmap <= 16'b0000111111110000;
		15'h2e46: char_row_bitmap <= 16'b0000111111110000;
		15'h2e47: char_row_bitmap <= 16'b0000000000000000;
		15'h2e48: char_row_bitmap <= 16'b0000000000000000;
		15'h2e49: char_row_bitmap <= 16'b0000111111110000;
		15'h2e4a: char_row_bitmap <= 16'b0000111111110000;
		15'h2e4b: char_row_bitmap <= 16'b0000000000000000;
		15'h2e4c: char_row_bitmap <= 16'b0000000000000000;
		15'h2e4d: char_row_bitmap <= 16'b0000111111110000;
		15'h2e4e: char_row_bitmap <= 16'b0000111111110000;
		15'h2e4f: char_row_bitmap <= 16'b0000000000000000;
		15'h2e50: char_row_bitmap <= 16'b0000000000000000;
		15'h2e51: char_row_bitmap <= 16'b0000000000000000;
		15'h2e52: char_row_bitmap <= 16'b0000000000000000;
		15'h2e53: char_row_bitmap <= 16'b0000000000000000;
		15'h2e54: char_row_bitmap <= 16'b0000000000000000;
		15'h2e55: char_row_bitmap <= 16'b0000000000000000;
		15'h2e56: char_row_bitmap <= 16'b0000000000000000;
		15'h2e57: char_row_bitmap <= 16'b0000000000000000;
		15'h2e58: char_row_bitmap <= 16'b0000000000000000;
		15'h2e59: char_row_bitmap <= 16'b0000011111100000;
		15'h2e5a: char_row_bitmap <= 16'b0000111111110000;
		15'h2e5b: char_row_bitmap <= 16'b0001110110111000;
		15'h2e5c: char_row_bitmap <= 16'b0001100000011000;
		15'h2e5d: char_row_bitmap <= 16'b0001110000111000;
		15'h2e5e: char_row_bitmap <= 16'b0001110000111000;
		15'h2e5f: char_row_bitmap <= 16'b0001100000011000;
		15'h2e60: char_row_bitmap <= 16'b0001110110111000;
		15'h2e61: char_row_bitmap <= 16'b0000111111110000;
		15'h2e62: char_row_bitmap <= 16'b0000011111100000;
		15'h2e63: char_row_bitmap <= 16'b0000000000000000;
		15'h2e64: char_row_bitmap <= 16'b0000000000000000;
		15'h2e65: char_row_bitmap <= 16'b0000000000000000;
		15'h2e66: char_row_bitmap <= 16'b0000000000000000;
		15'h2e67: char_row_bitmap <= 16'b0000000000000000;
		15'h2e68: char_row_bitmap <= 16'b0000000000000000;
		15'h2e69: char_row_bitmap <= 16'b0000000000000000;
		15'h2e6a: char_row_bitmap <= 16'b0000000000000000;
		15'h2e6b: char_row_bitmap <= 16'b0111111111111110;
		15'h2e6c: char_row_bitmap <= 16'b0111111111111110;
		15'h2e6d: char_row_bitmap <= 16'b0110000000000110;
		15'h2e6e: char_row_bitmap <= 16'b0110000110000110;
		15'h2e6f: char_row_bitmap <= 16'b0110000110000110;
		15'h2e70: char_row_bitmap <= 16'b0110000110000110;
		15'h2e71: char_row_bitmap <= 16'b0110111111110110;
		15'h2e72: char_row_bitmap <= 16'b0110111111110110;
		15'h2e73: char_row_bitmap <= 16'b0110000110000110;
		15'h2e74: char_row_bitmap <= 16'b0110000110000110;
		15'h2e75: char_row_bitmap <= 16'b0110000110000110;
		15'h2e76: char_row_bitmap <= 16'b0110000000000110;
		15'h2e77: char_row_bitmap <= 16'b0111111111111110;
		15'h2e78: char_row_bitmap <= 16'b0111111111111110;
		15'h2e79: char_row_bitmap <= 16'b0000000000000000;
		15'h2e7a: char_row_bitmap <= 16'b0000000000000000;
		15'h2e7b: char_row_bitmap <= 16'b0000000000000000;
		15'h2e7c: char_row_bitmap <= 16'b0000000000000000;
		15'h2e7d: char_row_bitmap <= 16'b0000000000000000;
		15'h2e7e: char_row_bitmap <= 16'b0000000000000000;
		15'h2e7f: char_row_bitmap <= 16'b0111111111111110;
		15'h2e80: char_row_bitmap <= 16'b0111111111111110;
		15'h2e81: char_row_bitmap <= 16'b0110000000000110;
		15'h2e82: char_row_bitmap <= 16'b0110000000000110;
		15'h2e83: char_row_bitmap <= 16'b0110000000000110;
		15'h2e84: char_row_bitmap <= 16'b0110000000000110;
		15'h2e85: char_row_bitmap <= 16'b0110111111110110;
		15'h2e86: char_row_bitmap <= 16'b0110111111110110;
		15'h2e87: char_row_bitmap <= 16'b0110000000000110;
		15'h2e88: char_row_bitmap <= 16'b0110000000000110;
		15'h2e89: char_row_bitmap <= 16'b0110000000000110;
		15'h2e8a: char_row_bitmap <= 16'b0110000000000110;
		15'h2e8b: char_row_bitmap <= 16'b0111111111111110;
		15'h2e8c: char_row_bitmap <= 16'b0111111111111110;
		15'h2e8d: char_row_bitmap <= 16'b0000000000000000;
		15'h2e8e: char_row_bitmap <= 16'b0000000000000000;
		15'h2e8f: char_row_bitmap <= 16'b0000000000000000;
		15'h2e90: char_row_bitmap <= 16'b0000000000000000;
		15'h2e91: char_row_bitmap <= 16'b0000000000000000;
		15'h2e92: char_row_bitmap <= 16'b0000000000000000;
		15'h2e93: char_row_bitmap <= 16'b0111111111100000;
		15'h2e94: char_row_bitmap <= 16'b0111111111100000;
		15'h2e95: char_row_bitmap <= 16'b0110000000000110;
		15'h2e96: char_row_bitmap <= 16'b0110000000001110;
		15'h2e97: char_row_bitmap <= 16'b0110000000011100;
		15'h2e98: char_row_bitmap <= 16'b0110110000111000;
		15'h2e99: char_row_bitmap <= 16'b0110111001110000;
		15'h2e9a: char_row_bitmap <= 16'b0110011111100000;
		15'h2e9b: char_row_bitmap <= 16'b0110001111000110;
		15'h2e9c: char_row_bitmap <= 16'b0110000110000110;
		15'h2e9d: char_row_bitmap <= 16'b0110000000000110;
		15'h2e9e: char_row_bitmap <= 16'b0110000000000110;
		15'h2e9f: char_row_bitmap <= 16'b0111111111111110;
		15'h2ea0: char_row_bitmap <= 16'b0111111111111110;
		15'h2ea1: char_row_bitmap <= 16'b0000000000000000;
		15'h2ea2: char_row_bitmap <= 16'b0000000000000000;
		15'h2ea3: char_row_bitmap <= 16'b0000000000000000;
		15'h2ea4: char_row_bitmap <= 16'b0000000000000000;
		15'h2ea5: char_row_bitmap <= 16'b0000000000000000;
		15'h2ea6: char_row_bitmap <= 16'b0000000000000000;
		15'h2ea7: char_row_bitmap <= 16'b0111111111111110;
		15'h2ea8: char_row_bitmap <= 16'b0111111111111110;
		15'h2ea9: char_row_bitmap <= 16'b0110000000000110;
		15'h2eaa: char_row_bitmap <= 16'b0110000000000110;
		15'h2eab: char_row_bitmap <= 16'b0110000000000110;
		15'h2eac: char_row_bitmap <= 16'b0110000000000110;
		15'h2ead: char_row_bitmap <= 16'b0110000000000110;
		15'h2eae: char_row_bitmap <= 16'b0110000000000110;
		15'h2eaf: char_row_bitmap <= 16'b0110000000000110;
		15'h2eb0: char_row_bitmap <= 16'b0110000000000110;
		15'h2eb1: char_row_bitmap <= 16'b0110000000000110;
		15'h2eb2: char_row_bitmap <= 16'b0110000000000110;
		15'h2eb3: char_row_bitmap <= 16'b0111111111111110;
		15'h2eb4: char_row_bitmap <= 16'b0111111111111110;
		15'h2eb5: char_row_bitmap <= 16'b0000000000000000;
		15'h2eb6: char_row_bitmap <= 16'b0000000000000000;
		15'h2eb7: char_row_bitmap <= 16'b0000000000000000;
		15'h2eb8: char_row_bitmap <= 16'b0000000000000000;
		15'h2eb9: char_row_bitmap <= 16'b0000000000000000;
		15'h2eba: char_row_bitmap <= 16'b0000000000000000;
		15'h2ebb: char_row_bitmap <= 16'b0111111111111110;
		15'h2ebc: char_row_bitmap <= 16'b0111111111111110;
		15'h2ebd: char_row_bitmap <= 16'b0110000000000110;
		15'h2ebe: char_row_bitmap <= 16'b0110110000110110;
		15'h2ebf: char_row_bitmap <= 16'b0110111001110110;
		15'h2ec0: char_row_bitmap <= 16'b0110011111100110;
		15'h2ec1: char_row_bitmap <= 16'b0110001111000110;
		15'h2ec2: char_row_bitmap <= 16'b0110001111000110;
		15'h2ec3: char_row_bitmap <= 16'b0110011111100110;
		15'h2ec4: char_row_bitmap <= 16'b0110111001110110;
		15'h2ec5: char_row_bitmap <= 16'b0110110000110110;
		15'h2ec6: char_row_bitmap <= 16'b0110000000000110;
		15'h2ec7: char_row_bitmap <= 16'b0111111111111110;
		15'h2ec8: char_row_bitmap <= 16'b0111111111111110;
		15'h2ec9: char_row_bitmap <= 16'b0000000000000000;
		15'h2eca: char_row_bitmap <= 16'b0000000000000000;
		15'h2ecb: char_row_bitmap <= 16'b0000000000000000;
		15'h2ecc: char_row_bitmap <= 16'b0000000000000000;
		15'h2ecd: char_row_bitmap <= 16'b0000000000000000;
		15'h2ece: char_row_bitmap <= 16'b0000000000000000;
		15'h2ecf: char_row_bitmap <= 16'b0000000000000000;
		15'h2ed0: char_row_bitmap <= 16'b0000000000000000;
		15'h2ed1: char_row_bitmap <= 16'b0001111111111000;
		15'h2ed2: char_row_bitmap <= 16'b0001111111111000;
		15'h2ed3: char_row_bitmap <= 16'b0001111001111000;
		15'h2ed4: char_row_bitmap <= 16'b0001111001111000;
		15'h2ed5: char_row_bitmap <= 16'b0001100000011000;
		15'h2ed6: char_row_bitmap <= 16'b0001100000011000;
		15'h2ed7: char_row_bitmap <= 16'b0001111001111000;
		15'h2ed8: char_row_bitmap <= 16'b0001111001111000;
		15'h2ed9: char_row_bitmap <= 16'b0001111111111000;
		15'h2eda: char_row_bitmap <= 16'b0001111111111000;
		15'h2edb: char_row_bitmap <= 16'b0000000000000000;
		15'h2edc: char_row_bitmap <= 16'b0000000000000000;
		15'h2edd: char_row_bitmap <= 16'b0000000000000000;
		15'h2ede: char_row_bitmap <= 16'b0000000000000000;
		15'h2edf: char_row_bitmap <= 16'b0000000000000000;
		15'h2ee0: char_row_bitmap <= 16'b0000000000000000;
		15'h2ee1: char_row_bitmap <= 16'b0000000000000000;
		15'h2ee2: char_row_bitmap <= 16'b0000000000000000;
		15'h2ee3: char_row_bitmap <= 16'b0000000000000000;
		15'h2ee4: char_row_bitmap <= 16'b0000000000000000;
		15'h2ee5: char_row_bitmap <= 16'b0001111111111000;
		15'h2ee6: char_row_bitmap <= 16'b0001111111111000;
		15'h2ee7: char_row_bitmap <= 16'b0001111111111000;
		15'h2ee8: char_row_bitmap <= 16'b0001111111111000;
		15'h2ee9: char_row_bitmap <= 16'b0001100000011000;
		15'h2eea: char_row_bitmap <= 16'b0001100000011000;
		15'h2eeb: char_row_bitmap <= 16'b0001111111111000;
		15'h2eec: char_row_bitmap <= 16'b0001111111111000;
		15'h2eed: char_row_bitmap <= 16'b0001111111111000;
		15'h2eee: char_row_bitmap <= 16'b0001111111111000;
		15'h2eef: char_row_bitmap <= 16'b0000000000000000;
		15'h2ef0: char_row_bitmap <= 16'b0000000000000000;
		15'h2ef1: char_row_bitmap <= 16'b0000000000000000;
		15'h2ef2: char_row_bitmap <= 16'b0000000000000000;
		15'h2ef3: char_row_bitmap <= 16'b0000000000000000;
		15'h2ef4: char_row_bitmap <= 16'b0000000000000000;
		15'h2ef5: char_row_bitmap <= 16'b0000000000000000;
		15'h2ef6: char_row_bitmap <= 16'b0000000000000000;
		15'h2ef7: char_row_bitmap <= 16'b0000000000000000;
		15'h2ef8: char_row_bitmap <= 16'b0000000000000000;
		15'h2ef9: char_row_bitmap <= 16'b0000011111100000;
		15'h2efa: char_row_bitmap <= 16'b0000111111110000;
		15'h2efb: char_row_bitmap <= 16'b0001111001111000;
		15'h2efc: char_row_bitmap <= 16'b0001111001111000;
		15'h2efd: char_row_bitmap <= 16'b0001100000011000;
		15'h2efe: char_row_bitmap <= 16'b0001100000011000;
		15'h2eff: char_row_bitmap <= 16'b0001111001111000;
		15'h2f00: char_row_bitmap <= 16'b0001111001111000;
		15'h2f01: char_row_bitmap <= 16'b0000111111110000;
		15'h2f02: char_row_bitmap <= 16'b0000011111100000;
		15'h2f03: char_row_bitmap <= 16'b0000000000000000;
		15'h2f04: char_row_bitmap <= 16'b0000000000000000;
		15'h2f05: char_row_bitmap <= 16'b0000000000000000;
		15'h2f06: char_row_bitmap <= 16'b0000000000000000;
		15'h2f07: char_row_bitmap <= 16'b0000000000000000;
		15'h2f08: char_row_bitmap <= 16'b0000000000000000;
		15'h2f09: char_row_bitmap <= 16'b0000000000000000;
		15'h2f0a: char_row_bitmap <= 16'b0000000000000000;
		15'h2f0b: char_row_bitmap <= 16'b0000000000000000;
		15'h2f0c: char_row_bitmap <= 16'b0000000000000000;
		15'h2f0d: char_row_bitmap <= 16'b0000011111100000;
		15'h2f0e: char_row_bitmap <= 16'b0000111111110000;
		15'h2f0f: char_row_bitmap <= 16'b0001111111111000;
		15'h2f10: char_row_bitmap <= 16'b0001111111111000;
		15'h2f11: char_row_bitmap <= 16'b0001100000011000;
		15'h2f12: char_row_bitmap <= 16'b0001100000011000;
		15'h2f13: char_row_bitmap <= 16'b0001111111111000;
		15'h2f14: char_row_bitmap <= 16'b0001111111111000;
		15'h2f15: char_row_bitmap <= 16'b0000111111110000;
		15'h2f16: char_row_bitmap <= 16'b0000011111100000;
		15'h2f17: char_row_bitmap <= 16'b0000000000000000;
		15'h2f18: char_row_bitmap <= 16'b0000000000000000;
		15'h2f19: char_row_bitmap <= 16'b0000000000000000;
		15'h2f1a: char_row_bitmap <= 16'b0000000000000000;
		15'h2f1b: char_row_bitmap <= 16'b0000000000000000;
		15'h2f1c: char_row_bitmap <= 16'b0000000000000000;
		15'h2f1d: char_row_bitmap <= 16'b0000000000000000;
		15'h2f1e: char_row_bitmap <= 16'b0000000000000000;
		15'h2f1f: char_row_bitmap <= 16'b0000011111100000;
		15'h2f20: char_row_bitmap <= 16'b0000111111110000;
		15'h2f21: char_row_bitmap <= 16'b0001110000111000;
		15'h2f22: char_row_bitmap <= 16'b0011100000011100;
		15'h2f23: char_row_bitmap <= 16'b0111000110001110;
		15'h2f24: char_row_bitmap <= 16'b0110000110000110;
		15'h2f25: char_row_bitmap <= 16'b0110011111100110;
		15'h2f26: char_row_bitmap <= 16'b0110011111100110;
		15'h2f27: char_row_bitmap <= 16'b0110000110000110;
		15'h2f28: char_row_bitmap <= 16'b0111000110001110;
		15'h2f29: char_row_bitmap <= 16'b0011100000011100;
		15'h2f2a: char_row_bitmap <= 16'b0001110000111000;
		15'h2f2b: char_row_bitmap <= 16'b0000111111110000;
		15'h2f2c: char_row_bitmap <= 16'b0000011111100000;
		15'h2f2d: char_row_bitmap <= 16'b0000000000000000;
		15'h2f2e: char_row_bitmap <= 16'b0000000000000000;
		15'h2f2f: char_row_bitmap <= 16'b0000000000000000;
		15'h2f30: char_row_bitmap <= 16'b0000000000000000;
		15'h2f31: char_row_bitmap <= 16'b0000000000000000;
		15'h2f32: char_row_bitmap <= 16'b0000000000000000;
		15'h2f33: char_row_bitmap <= 16'b0000011111100000;
		15'h2f34: char_row_bitmap <= 16'b0000111111110000;
		15'h2f35: char_row_bitmap <= 16'b0001110000111000;
		15'h2f36: char_row_bitmap <= 16'b0011100000011100;
		15'h2f37: char_row_bitmap <= 16'b0111000000001110;
		15'h2f38: char_row_bitmap <= 16'b0110000000000110;
		15'h2f39: char_row_bitmap <= 16'b0110000000000110;
		15'h2f3a: char_row_bitmap <= 16'b0110000000000110;
		15'h2f3b: char_row_bitmap <= 16'b0110000000000110;
		15'h2f3c: char_row_bitmap <= 16'b0111000000001110;
		15'h2f3d: char_row_bitmap <= 16'b0011100000011100;
		15'h2f3e: char_row_bitmap <= 16'b0001110000111000;
		15'h2f3f: char_row_bitmap <= 16'b0000111111110000;
		15'h2f40: char_row_bitmap <= 16'b0000011111100000;
		15'h2f41: char_row_bitmap <= 16'b0000000000000000;
		15'h2f42: char_row_bitmap <= 16'b0000000000000000;
		15'h2f43: char_row_bitmap <= 16'b0000000000000000;
		15'h2f44: char_row_bitmap <= 16'b0000000000000000;
		15'h2f45: char_row_bitmap <= 16'b0000000000000000;
		15'h2f46: char_row_bitmap <= 16'b0000000000000000;
		15'h2f47: char_row_bitmap <= 16'b0000011111100000;
		15'h2f48: char_row_bitmap <= 16'b0000111111110000;
		15'h2f49: char_row_bitmap <= 16'b0001110000111000;
		15'h2f4a: char_row_bitmap <= 16'b0011100000011100;
		15'h2f4b: char_row_bitmap <= 16'b0111001111001110;
		15'h2f4c: char_row_bitmap <= 16'b0110011111100110;
		15'h2f4d: char_row_bitmap <= 16'b0110011111100110;
		15'h2f4e: char_row_bitmap <= 16'b0110011111100110;
		15'h2f4f: char_row_bitmap <= 16'b0110011111100110;
		15'h2f50: char_row_bitmap <= 16'b0111001111001110;
		15'h2f51: char_row_bitmap <= 16'b0011100000011100;
		15'h2f52: char_row_bitmap <= 16'b0001110000111000;
		15'h2f53: char_row_bitmap <= 16'b0000111111110000;
		15'h2f54: char_row_bitmap <= 16'b0000011111100000;
		15'h2f55: char_row_bitmap <= 16'b0000000000000000;
		15'h2f56: char_row_bitmap <= 16'b0000000000000000;
		15'h2f57: char_row_bitmap <= 16'b0000000000000000;
		15'h2f58: char_row_bitmap <= 16'b0000000000000000;
		15'h2f59: char_row_bitmap <= 16'b0000000000000000;
		15'h2f5a: char_row_bitmap <= 16'b0000000000001100;
		15'h2f5b: char_row_bitmap <= 16'b0000000000001100;
		15'h2f5c: char_row_bitmap <= 16'b0000000000011100;
		15'h2f5d: char_row_bitmap <= 16'b0000000000011000;
		15'h2f5e: char_row_bitmap <= 16'b0000000000111000;
		15'h2f5f: char_row_bitmap <= 16'b0000000011110000;
		15'h2f60: char_row_bitmap <= 16'b1100000111100000;
		15'h2f61: char_row_bitmap <= 16'b1110000110000000;
		15'h2f62: char_row_bitmap <= 16'b0111001100000000;
		15'h2f63: char_row_bitmap <= 16'b0011001100000000;
		15'h2f64: char_row_bitmap <= 16'b0001111000000000;
		15'h2f65: char_row_bitmap <= 16'b0001111000000000;
		15'h2f66: char_row_bitmap <= 16'b0000110000000000;
		15'h2f67: char_row_bitmap <= 16'b0000110000000000;
		15'h2f68: char_row_bitmap <= 16'b0000000000000000;
		15'h2f69: char_row_bitmap <= 16'b0000000000000000;
		15'h2f6a: char_row_bitmap <= 16'b0000000000000000;
		15'h2f6b: char_row_bitmap <= 16'b0000000000000000;
		15'h2f6c: char_row_bitmap <= 16'b0000000000000000;
		15'h2f6d: char_row_bitmap <= 16'b0000000000000000;
		15'h2f6e: char_row_bitmap <= 16'b0000000000000000;
		15'h2f6f: char_row_bitmap <= 16'b0000000000000000;
		15'h2f70: char_row_bitmap <= 16'b0000110000000000;
		15'h2f71: char_row_bitmap <= 16'b0000110000000000;
		15'h2f72: char_row_bitmap <= 16'b0001111000000000;
		15'h2f73: char_row_bitmap <= 16'b0001111000000000;
		15'h2f74: char_row_bitmap <= 16'b0011001100000000;
		15'h2f75: char_row_bitmap <= 16'b0111001100000000;
		15'h2f76: char_row_bitmap <= 16'b1110000110000000;
		15'h2f77: char_row_bitmap <= 16'b1100000111100000;
		15'h2f78: char_row_bitmap <= 16'b0000000011110000;
		15'h2f79: char_row_bitmap <= 16'b0000000000111000;
		15'h2f7a: char_row_bitmap <= 16'b0000000000011000;
		15'h2f7b: char_row_bitmap <= 16'b0000000000011100;
		15'h2f7c: char_row_bitmap <= 16'b0000000000001100;
		15'h2f7d: char_row_bitmap <= 16'b0000000000001100;
		15'h2f7e: char_row_bitmap <= 16'b0000000000000000;
		15'h2f7f: char_row_bitmap <= 16'b0000000000000000;
		15'h2f80: char_row_bitmap <= 16'b0000000000000000;
		15'h2f81: char_row_bitmap <= 16'b0000000000000000;
		15'h2f82: char_row_bitmap <= 16'b0000000000000000;
		15'h2f83: char_row_bitmap <= 16'b0000000000000000;
		15'h2f84: char_row_bitmap <= 16'b0000000000000000;
		15'h2f85: char_row_bitmap <= 16'b0000000000000000;
		15'h2f86: char_row_bitmap <= 16'b0000000000000000;
		15'h2f87: char_row_bitmap <= 16'b0000000000000000;
		15'h2f88: char_row_bitmap <= 16'b0000000000000000;
		15'h2f89: char_row_bitmap <= 16'b0000000000000000;
		15'h2f8a: char_row_bitmap <= 16'b0000011111111111;
		15'h2f8b: char_row_bitmap <= 16'b0001111111111111;
		15'h2f8c: char_row_bitmap <= 16'b0011110000000000;
		15'h2f8d: char_row_bitmap <= 16'b0111000000000000;
		15'h2f8e: char_row_bitmap <= 16'b0110000000000000;
		15'h2f8f: char_row_bitmap <= 16'b1110000000000000;
		15'h2f90: char_row_bitmap <= 16'b1100000000000000;
		15'h2f91: char_row_bitmap <= 16'b1100000000000000;
		15'h2f92: char_row_bitmap <= 16'b0000000000000000;
		15'h2f93: char_row_bitmap <= 16'b0000000000000000;
		15'h2f94: char_row_bitmap <= 16'b0000000000000000;
		15'h2f95: char_row_bitmap <= 16'b0000000000000000;
		15'h2f96: char_row_bitmap <= 16'b0000000000000000;
		15'h2f97: char_row_bitmap <= 16'b0000000000000000;
		15'h2f98: char_row_bitmap <= 16'b0000000000000000;
		15'h2f99: char_row_bitmap <= 16'b0000000000000000;
		15'h2f9a: char_row_bitmap <= 16'b0000000000000000;
		15'h2f9b: char_row_bitmap <= 16'b0000000000000000;
		15'h2f9c: char_row_bitmap <= 16'b0000000000000000;
		15'h2f9d: char_row_bitmap <= 16'b0000000000000000;
		15'h2f9e: char_row_bitmap <= 16'b1111111110000000;
		15'h2f9f: char_row_bitmap <= 16'b1111111111100000;
		15'h2fa0: char_row_bitmap <= 16'b0000000011110000;
		15'h2fa1: char_row_bitmap <= 16'b0000000000111000;
		15'h2fa2: char_row_bitmap <= 16'b0000000000011000;
		15'h2fa3: char_row_bitmap <= 16'b0000000000011100;
		15'h2fa4: char_row_bitmap <= 16'b0000000000001100;
		15'h2fa5: char_row_bitmap <= 16'b0000000000001100;
		15'h2fa6: char_row_bitmap <= 16'b0000000000000000;
		15'h2fa7: char_row_bitmap <= 16'b0000000000000000;
		15'h2fa8: char_row_bitmap <= 16'b0000000000000000;
		15'h2fa9: char_row_bitmap <= 16'b0000000000000000;
		15'h2faa: char_row_bitmap <= 16'b0000000000000000;
		15'h2fab: char_row_bitmap <= 16'b0000000000000000;
		15'h2fac: char_row_bitmap <= 16'b0000001100000000;
		15'h2fad: char_row_bitmap <= 16'b0000001100000000;
		15'h2fae: char_row_bitmap <= 16'b0000011110000000;
		15'h2faf: char_row_bitmap <= 16'b0000011110000000;
		15'h2fb0: char_row_bitmap <= 16'b0000110011000000;
		15'h2fb1: char_row_bitmap <= 16'b0001110011100000;
		15'h2fb2: char_row_bitmap <= 16'b1111100001111111;
		15'h2fb3: char_row_bitmap <= 16'b1111000000111111;
		15'h2fb4: char_row_bitmap <= 16'b0000000000000000;
		15'h2fb5: char_row_bitmap <= 16'b0000000000000000;
		15'h2fb6: char_row_bitmap <= 16'b0000000000000000;
		15'h2fb7: char_row_bitmap <= 16'b0000000000000000;
		15'h2fb8: char_row_bitmap <= 16'b0000000000000000;
		15'h2fb9: char_row_bitmap <= 16'b0000000000000000;
		15'h2fba: char_row_bitmap <= 16'b0000000000000000;
		15'h2fbb: char_row_bitmap <= 16'b0000000000000000;
		15'h2fbc: char_row_bitmap <= 16'b0000000000000000;
		15'h2fbd: char_row_bitmap <= 16'b0000000000000000;
		15'h2fbe: char_row_bitmap <= 16'b0000000000000000;
		15'h2fbf: char_row_bitmap <= 16'b0000000000000000;
		15'h2fc0: char_row_bitmap <= 16'b0000000000000011;
		15'h2fc1: char_row_bitmap <= 16'b0000000000000011;
		15'h2fc2: char_row_bitmap <= 16'b0000000000000111;
		15'h2fc3: char_row_bitmap <= 16'b0000000000000111;
		15'h2fc4: char_row_bitmap <= 16'b0000000000001100;
		15'h2fc5: char_row_bitmap <= 16'b0000000000111100;
		15'h2fc6: char_row_bitmap <= 16'b0000011111111000;
		15'h2fc7: char_row_bitmap <= 16'b0001111111100000;
		15'h2fc8: char_row_bitmap <= 16'b0011110000000000;
		15'h2fc9: char_row_bitmap <= 16'b0111000000000000;
		15'h2fca: char_row_bitmap <= 16'b0110000000000000;
		15'h2fcb: char_row_bitmap <= 16'b1110000000000000;
		15'h2fcc: char_row_bitmap <= 16'b1100000000000000;
		15'h2fcd: char_row_bitmap <= 16'b1100000000000000;
		15'h2fce: char_row_bitmap <= 16'b0000000000000000;
		15'h2fcf: char_row_bitmap <= 16'b0000000000000000;
		15'h2fd0: char_row_bitmap <= 16'b0000000000000000;
		15'h2fd1: char_row_bitmap <= 16'b0000000000000000;
		15'h2fd2: char_row_bitmap <= 16'b0000000000000000;
		15'h2fd3: char_row_bitmap <= 16'b0000000000000000;
		15'h2fd4: char_row_bitmap <= 16'b0000000000000000;
		15'h2fd5: char_row_bitmap <= 16'b0000000000000000;
		15'h2fd6: char_row_bitmap <= 16'b1000000000000000;
		15'h2fd7: char_row_bitmap <= 16'b1000000000000000;
		15'h2fd8: char_row_bitmap <= 16'b1100000000000000;
		15'h2fd9: char_row_bitmap <= 16'b1110000000000000;
		15'h2fda: char_row_bitmap <= 16'b0111111110000000;
		15'h2fdb: char_row_bitmap <= 16'b0011111111100000;
		15'h2fdc: char_row_bitmap <= 16'b0000000011110000;
		15'h2fdd: char_row_bitmap <= 16'b0000000000111000;
		15'h2fde: char_row_bitmap <= 16'b0000000000011000;
		15'h2fdf: char_row_bitmap <= 16'b0000000000011100;
		15'h2fe0: char_row_bitmap <= 16'b0000000000001100;
		15'h2fe1: char_row_bitmap <= 16'b0000000000001100;
		15'h2fe2: char_row_bitmap <= 16'b0000000000000000;
		15'h2fe3: char_row_bitmap <= 16'b0000000000000000;
		15'h2fe4: char_row_bitmap <= 16'b0000000000000000;
		15'h2fe5: char_row_bitmap <= 16'b0000000000000000;
		15'h2fe6: char_row_bitmap <= 16'b0000000000000000;
		15'h2fe7: char_row_bitmap <= 16'b0000000000000000;
		15'h2fe8: char_row_bitmap <= 16'b0000000000000011;
		15'h2fe9: char_row_bitmap <= 16'b0000000000000011;
		15'h2fea: char_row_bitmap <= 16'b0000000000000111;
		15'h2feb: char_row_bitmap <= 16'b0000000000000111;
		15'h2fec: char_row_bitmap <= 16'b0000000000001100;
		15'h2fed: char_row_bitmap <= 16'b0000000000111100;
		15'h2fee: char_row_bitmap <= 16'b1111111111111000;
		15'h2fef: char_row_bitmap <= 16'b1111111111110000;
		15'h2ff0: char_row_bitmap <= 16'b0000000000000000;
		15'h2ff1: char_row_bitmap <= 16'b0000000000000000;
		15'h2ff2: char_row_bitmap <= 16'b0000000000000000;
		15'h2ff3: char_row_bitmap <= 16'b0000000000000000;
		15'h2ff4: char_row_bitmap <= 16'b0000000000000000;
		15'h2ff5: char_row_bitmap <= 16'b0000000000000000;
		15'h2ff6: char_row_bitmap <= 16'b0000000000000000;
		15'h2ff7: char_row_bitmap <= 16'b0000000000000000;
		15'h2ff8: char_row_bitmap <= 16'b0000000000000000;
		15'h2ff9: char_row_bitmap <= 16'b0000000000000000;
		15'h2ffa: char_row_bitmap <= 16'b0000000000000000;
		15'h2ffb: char_row_bitmap <= 16'b0000000000000000;
		15'h2ffc: char_row_bitmap <= 16'b0000000000000000;
		15'h2ffd: char_row_bitmap <= 16'b0000000000000000;
		15'h2ffe: char_row_bitmap <= 16'b1000000000000000;
		15'h2fff: char_row_bitmap <= 16'b1000000000000000;
		15'h3000: char_row_bitmap <= 16'b1100000000000000;
		15'h3001: char_row_bitmap <= 16'b1110000000000000;
		15'h3002: char_row_bitmap <= 16'b0111111111111111;
		15'h3003: char_row_bitmap <= 16'b0011111111111111;
		15'h3004: char_row_bitmap <= 16'b0000000000000000;
		15'h3005: char_row_bitmap <= 16'b0000000000000000;
		15'h3006: char_row_bitmap <= 16'b0000000000000000;
		15'h3007: char_row_bitmap <= 16'b0000000000000000;
		15'h3008: char_row_bitmap <= 16'b0000000000000000;
		15'h3009: char_row_bitmap <= 16'b0000000000000000;
		15'h300a: char_row_bitmap <= 16'b0000000000000000;
		15'h300b: char_row_bitmap <= 16'b0000000000000000;
		15'h300c: char_row_bitmap <= 16'b0000000000000000;
		15'h300d: char_row_bitmap <= 16'b0000000000000000;
		15'h300e: char_row_bitmap <= 16'b1100000000000000;
		15'h300f: char_row_bitmap <= 16'b1100000000000000;
		15'h3010: char_row_bitmap <= 16'b1110000000000000;
		15'h3011: char_row_bitmap <= 16'b0110000000000000;
		15'h3012: char_row_bitmap <= 16'b0111000000000000;
		15'h3013: char_row_bitmap <= 16'b0011110000000000;
		15'h3014: char_row_bitmap <= 16'b0001111111111111;
		15'h3015: char_row_bitmap <= 16'b0000011111111111;
		15'h3016: char_row_bitmap <= 16'b0000000000000000;
		15'h3017: char_row_bitmap <= 16'b0000000000000000;
		15'h3018: char_row_bitmap <= 16'b0000000000000000;
		15'h3019: char_row_bitmap <= 16'b0000000000000000;
		15'h301a: char_row_bitmap <= 16'b0000000000000000;
		15'h301b: char_row_bitmap <= 16'b0000000000000000;
		15'h301c: char_row_bitmap <= 16'b0000000000000000;
		15'h301d: char_row_bitmap <= 16'b0000000000000000;
		15'h301e: char_row_bitmap <= 16'b0000000000000000;
		15'h301f: char_row_bitmap <= 16'b0000000000000000;
		15'h3020: char_row_bitmap <= 16'b0000000000000000;
		15'h3021: char_row_bitmap <= 16'b0000000000000000;
		15'h3022: char_row_bitmap <= 16'b0000000000001100;
		15'h3023: char_row_bitmap <= 16'b0000000000001100;
		15'h3024: char_row_bitmap <= 16'b0000000000011100;
		15'h3025: char_row_bitmap <= 16'b0000000000011000;
		15'h3026: char_row_bitmap <= 16'b0000000000111000;
		15'h3027: char_row_bitmap <= 16'b0000000011110000;
		15'h3028: char_row_bitmap <= 16'b1111111111100000;
		15'h3029: char_row_bitmap <= 16'b1111111110000000;
		15'h302a: char_row_bitmap <= 16'b0000000000000000;
		15'h302b: char_row_bitmap <= 16'b0000000000000000;
		15'h302c: char_row_bitmap <= 16'b0000000000000000;
		15'h302d: char_row_bitmap <= 16'b0000000000000000;
		15'h302e: char_row_bitmap <= 16'b0000000000000000;
		15'h302f: char_row_bitmap <= 16'b0000000000000000;
		15'h3030: char_row_bitmap <= 16'b0000000000000000;
		15'h3031: char_row_bitmap <= 16'b0000000000000000;
		15'h3032: char_row_bitmap <= 16'b0000000000000000;
		15'h3033: char_row_bitmap <= 16'b0000000000000000;
		15'h3034: char_row_bitmap <= 16'b0000000000000000;
		15'h3035: char_row_bitmap <= 16'b0000000000000000;
		15'h3036: char_row_bitmap <= 16'b0000000000000000;
		15'h3037: char_row_bitmap <= 16'b0000000000000000;
		15'h3038: char_row_bitmap <= 16'b0000000000000000;
		15'h3039: char_row_bitmap <= 16'b0000000000000000;
		15'h303a: char_row_bitmap <= 16'b0000000000000000;
		15'h303b: char_row_bitmap <= 16'b0000000000000000;
		15'h303c: char_row_bitmap <= 16'b1111000000111111;
		15'h303d: char_row_bitmap <= 16'b1111100001111111;
		15'h303e: char_row_bitmap <= 16'b0001110011100000;
		15'h303f: char_row_bitmap <= 16'b0000110011000000;
		15'h3040: char_row_bitmap <= 16'b0000011110000000;
		15'h3041: char_row_bitmap <= 16'b0000011110000000;
		15'h3042: char_row_bitmap <= 16'b0000001100000000;
		15'h3043: char_row_bitmap <= 16'b0000001100000000;
		15'h3044: char_row_bitmap <= 16'b0000000000000000;
		15'h3045: char_row_bitmap <= 16'b0000000000000000;
		15'h3046: char_row_bitmap <= 16'b0000000000000000;
		15'h3047: char_row_bitmap <= 16'b0000000000000000;
		15'h3048: char_row_bitmap <= 16'b0000000000000000;
		15'h3049: char_row_bitmap <= 16'b0000000000000000;
		15'h304a: char_row_bitmap <= 16'b1100000000000000;
		15'h304b: char_row_bitmap <= 16'b1100000000000000;
		15'h304c: char_row_bitmap <= 16'b1110000000000000;
		15'h304d: char_row_bitmap <= 16'b0110000000000000;
		15'h304e: char_row_bitmap <= 16'b0111000000000000;
		15'h304f: char_row_bitmap <= 16'b0011110000000000;
		15'h3050: char_row_bitmap <= 16'b0001111111100000;
		15'h3051: char_row_bitmap <= 16'b0000011111111000;
		15'h3052: char_row_bitmap <= 16'b0000000000111100;
		15'h3053: char_row_bitmap <= 16'b0000000000001100;
		15'h3054: char_row_bitmap <= 16'b0000000000000111;
		15'h3055: char_row_bitmap <= 16'b0000000000000111;
		15'h3056: char_row_bitmap <= 16'b0000000000000011;
		15'h3057: char_row_bitmap <= 16'b0000000000000011;
		15'h3058: char_row_bitmap <= 16'b0000000000000000;
		15'h3059: char_row_bitmap <= 16'b0000000000000000;
		15'h305a: char_row_bitmap <= 16'b0000000000000000;
		15'h305b: char_row_bitmap <= 16'b0000000000000000;
		15'h305c: char_row_bitmap <= 16'b0000000000000000;
		15'h305d: char_row_bitmap <= 16'b0000000000000000;
		15'h305e: char_row_bitmap <= 16'b0000000000001100;
		15'h305f: char_row_bitmap <= 16'b0000000000001100;
		15'h3060: char_row_bitmap <= 16'b0000000000011100;
		15'h3061: char_row_bitmap <= 16'b0000000000011000;
		15'h3062: char_row_bitmap <= 16'b0000000000111000;
		15'h3063: char_row_bitmap <= 16'b0000000011110000;
		15'h3064: char_row_bitmap <= 16'b0011111111100000;
		15'h3065: char_row_bitmap <= 16'b0111111110000000;
		15'h3066: char_row_bitmap <= 16'b1110000000000000;
		15'h3067: char_row_bitmap <= 16'b1100000000000000;
		15'h3068: char_row_bitmap <= 16'b1000000000000000;
		15'h3069: char_row_bitmap <= 16'b1000000000000000;
		15'h306a: char_row_bitmap <= 16'b0000000000000000;
		15'h306b: char_row_bitmap <= 16'b0000000000000000;
		15'h306c: char_row_bitmap <= 16'b0000000000000000;
		15'h306d: char_row_bitmap <= 16'b0000000000000000;
		15'h306e: char_row_bitmap <= 16'b0000000000000000;
		15'h306f: char_row_bitmap <= 16'b0000000000000000;
		15'h3070: char_row_bitmap <= 16'b0000000000000000;
		15'h3071: char_row_bitmap <= 16'b0000000000000000;
		15'h3072: char_row_bitmap <= 16'b0000000000000000;
		15'h3073: char_row_bitmap <= 16'b0000000000000000;
		15'h3074: char_row_bitmap <= 16'b0000000000000000;
		15'h3075: char_row_bitmap <= 16'b0000000000000000;
		15'h3076: char_row_bitmap <= 16'b0000000000000000;
		15'h3077: char_row_bitmap <= 16'b0000000000000000;
		15'h3078: char_row_bitmap <= 16'b1111111111110000;
		15'h3079: char_row_bitmap <= 16'b1111111111111000;
		15'h307a: char_row_bitmap <= 16'b0000000000111100;
		15'h307b: char_row_bitmap <= 16'b0000000000001100;
		15'h307c: char_row_bitmap <= 16'b0000000000000111;
		15'h307d: char_row_bitmap <= 16'b0000000000000111;
		15'h307e: char_row_bitmap <= 16'b0000000000000011;
		15'h307f: char_row_bitmap <= 16'b0000000000000011;
		15'h3080: char_row_bitmap <= 16'b0000000000000000;
		15'h3081: char_row_bitmap <= 16'b0000000000000000;
		15'h3082: char_row_bitmap <= 16'b0000000000000000;
		15'h3083: char_row_bitmap <= 16'b0000000000000000;
		15'h3084: char_row_bitmap <= 16'b0000000000000000;
		15'h3085: char_row_bitmap <= 16'b0000000000000000;
		15'h3086: char_row_bitmap <= 16'b0000000000000000;
		15'h3087: char_row_bitmap <= 16'b0000000000000000;
		15'h3088: char_row_bitmap <= 16'b0000000000000000;
		15'h3089: char_row_bitmap <= 16'b0000000000000000;
		15'h308a: char_row_bitmap <= 16'b0000000000000000;
		15'h308b: char_row_bitmap <= 16'b0000000000000000;
		15'h308c: char_row_bitmap <= 16'b0011111111111111;
		15'h308d: char_row_bitmap <= 16'b0111111111111111;
		15'h308e: char_row_bitmap <= 16'b1110000000000000;
		15'h308f: char_row_bitmap <= 16'b1100000000000000;
		15'h3090: char_row_bitmap <= 16'b1000000000000000;
		15'h3091: char_row_bitmap <= 16'b1000000000000000;
		15'h3092: char_row_bitmap <= 16'b0000000000000000;
		15'h3093: char_row_bitmap <= 16'b0000000000000000;
		15'h3094: char_row_bitmap <= 16'b0000000000000000;
		15'h3095: char_row_bitmap <= 16'b0000000000000000;
		15'h3096: char_row_bitmap <= 16'b0000000000000000;
		15'h3097: char_row_bitmap <= 16'b0000000000000000;
		15'h3098: char_row_bitmap <= 16'b0011100000000000;
		15'h3099: char_row_bitmap <= 16'b0011110000000000;
		15'h309a: char_row_bitmap <= 16'b0000111000000000;
		15'h309b: char_row_bitmap <= 16'b0000011000000000;
		15'h309c: char_row_bitmap <= 16'b0000011100000000;
		15'h309d: char_row_bitmap <= 16'b0000001110000000;
		15'h309e: char_row_bitmap <= 16'b0000000110000000;
		15'h309f: char_row_bitmap <= 16'b0000000110000000;
		15'h30a0: char_row_bitmap <= 16'b0000000111000000;
		15'h30a1: char_row_bitmap <= 16'b0000000011110000;
		15'h30a2: char_row_bitmap <= 16'b0000000000111100;
		15'h30a3: char_row_bitmap <= 16'b0000000000111100;
		15'h30a4: char_row_bitmap <= 16'b0000000011110000;
		15'h30a5: char_row_bitmap <= 16'b0000000111000000;
		15'h30a6: char_row_bitmap <= 16'b0000001110000000;
		15'h30a7: char_row_bitmap <= 16'b0000001100000000;
		15'h30a8: char_row_bitmap <= 16'b0000001100000000;
		15'h30a9: char_row_bitmap <= 16'b0000001100000000;
		15'h30aa: char_row_bitmap <= 16'b0000001100000000;
		15'h30ab: char_row_bitmap <= 16'b0000001100000000;
		15'h30ac: char_row_bitmap <= 16'b0000000000011100;
		15'h30ad: char_row_bitmap <= 16'b0000000000111100;
		15'h30ae: char_row_bitmap <= 16'b0000000001110000;
		15'h30af: char_row_bitmap <= 16'b0000000001100000;
		15'h30b0: char_row_bitmap <= 16'b0000000011100000;
		15'h30b1: char_row_bitmap <= 16'b0000000111000000;
		15'h30b2: char_row_bitmap <= 16'b0000000110000000;
		15'h30b3: char_row_bitmap <= 16'b0000000110000000;
		15'h30b4: char_row_bitmap <= 16'b0000001110000000;
		15'h30b5: char_row_bitmap <= 16'b0000111100000000;
		15'h30b6: char_row_bitmap <= 16'b0011110000000000;
		15'h30b7: char_row_bitmap <= 16'b0011110000000000;
		15'h30b8: char_row_bitmap <= 16'b0000111100000000;
		15'h30b9: char_row_bitmap <= 16'b0000001110000000;
		15'h30ba: char_row_bitmap <= 16'b0000000111000000;
		15'h30bb: char_row_bitmap <= 16'b0000000011000000;
		15'h30bc: char_row_bitmap <= 16'b0000000011000000;
		15'h30bd: char_row_bitmap <= 16'b0000000011000000;
		15'h30be: char_row_bitmap <= 16'b0000000011000000;
		15'h30bf: char_row_bitmap <= 16'b0000000011000000;
		15'h30c0: char_row_bitmap <= 16'b0011100000000000;
		15'h30c1: char_row_bitmap <= 16'b0011110000000000;
		15'h30c2: char_row_bitmap <= 16'b0000111000000000;
		15'h30c3: char_row_bitmap <= 16'b0000011000000000;
		15'h30c4: char_row_bitmap <= 16'b0000011100000000;
		15'h30c5: char_row_bitmap <= 16'b0000001100000000;
		15'h30c6: char_row_bitmap <= 16'b0000001100000000;
		15'h30c7: char_row_bitmap <= 16'b0000001100000000;
		15'h30c8: char_row_bitmap <= 16'b0000001100000000;
		15'h30c9: char_row_bitmap <= 16'b0000001100000000;
		15'h30ca: char_row_bitmap <= 16'b0000001100000000;
		15'h30cb: char_row_bitmap <= 16'b0000001100000000;
		15'h30cc: char_row_bitmap <= 16'b0000001100000000;
		15'h30cd: char_row_bitmap <= 16'b0000001100000000;
		15'h30ce: char_row_bitmap <= 16'b0000001100000000;
		15'h30cf: char_row_bitmap <= 16'b0000001100000000;
		15'h30d0: char_row_bitmap <= 16'b0000001100000000;
		15'h30d1: char_row_bitmap <= 16'b0000001100000000;
		15'h30d2: char_row_bitmap <= 16'b0000001100000000;
		15'h30d3: char_row_bitmap <= 16'b0000001100000000;
		15'h30d4: char_row_bitmap <= 16'b0000001100000000;
		15'h30d5: char_row_bitmap <= 16'b0000001100000000;
		15'h30d6: char_row_bitmap <= 16'b0000001100000000;
		15'h30d7: char_row_bitmap <= 16'b0000001100000000;
		15'h30d8: char_row_bitmap <= 16'b0000001100000000;
		15'h30d9: char_row_bitmap <= 16'b0000001100000000;
		15'h30da: char_row_bitmap <= 16'b0000001100000000;
		15'h30db: char_row_bitmap <= 16'b0000001100000000;
		15'h30dc: char_row_bitmap <= 16'b0000001100000000;
		15'h30dd: char_row_bitmap <= 16'b0000001100000000;
		15'h30de: char_row_bitmap <= 16'b0000001100000000;
		15'h30df: char_row_bitmap <= 16'b0000001100000000;
		15'h30e0: char_row_bitmap <= 16'b0000001100000000;
		15'h30e1: char_row_bitmap <= 16'b0000011100000000;
		15'h30e2: char_row_bitmap <= 16'b0000011000000000;
		15'h30e3: char_row_bitmap <= 16'b0000111000000000;
		15'h30e4: char_row_bitmap <= 16'b0011110000000000;
		15'h30e5: char_row_bitmap <= 16'b0011100000000000;
		15'h30e6: char_row_bitmap <= 16'b0000000000000000;
		15'h30e7: char_row_bitmap <= 16'b0000000000000000;
		15'h30e8: char_row_bitmap <= 16'b0000001100000000;
		15'h30e9: char_row_bitmap <= 16'b0000001100000000;
		15'h30ea: char_row_bitmap <= 16'b0000001100000000;
		15'h30eb: char_row_bitmap <= 16'b0000001100000000;
		15'h30ec: char_row_bitmap <= 16'b0000001100000000;
		15'h30ed: char_row_bitmap <= 16'b0000001110000000;
		15'h30ee: char_row_bitmap <= 16'b0000000111000000;
		15'h30ef: char_row_bitmap <= 16'b0000000011110000;
		15'h30f0: char_row_bitmap <= 16'b0000000000111100;
		15'h30f1: char_row_bitmap <= 16'b0000000000111100;
		15'h30f2: char_row_bitmap <= 16'b0000000011110000;
		15'h30f3: char_row_bitmap <= 16'b0000000111000000;
		15'h30f4: char_row_bitmap <= 16'b0000001110000000;
		15'h30f5: char_row_bitmap <= 16'b0000001100000000;
		15'h30f6: char_row_bitmap <= 16'b0000001100000000;
		15'h30f7: char_row_bitmap <= 16'b0000001100000000;
		15'h30f8: char_row_bitmap <= 16'b0000001100000000;
		15'h30f9: char_row_bitmap <= 16'b0000001100000000;
		15'h30fa: char_row_bitmap <= 16'b0000001100000000;
		15'h30fb: char_row_bitmap <= 16'b0000001100000000;
		15'h30fc: char_row_bitmap <= 16'b0011100000000000;
		15'h30fd: char_row_bitmap <= 16'b0011110000000000;
		15'h30fe: char_row_bitmap <= 16'b0000111000000000;
		15'h30ff: char_row_bitmap <= 16'b0000011000000000;
		15'h3100: char_row_bitmap <= 16'b0000011100000000;
		15'h3101: char_row_bitmap <= 16'b0000001100000000;
		15'h3102: char_row_bitmap <= 16'b0000001100000000;
		15'h3103: char_row_bitmap <= 16'b0000001100000000;
		15'h3104: char_row_bitmap <= 16'b0000001100000000;
		15'h3105: char_row_bitmap <= 16'b0000001100000000;
		15'h3106: char_row_bitmap <= 16'b0000001100000000;
		15'h3107: char_row_bitmap <= 16'b0000001100000000;
		15'h3108: char_row_bitmap <= 16'b0000001100000000;
		15'h3109: char_row_bitmap <= 16'b0000001100000000;
		15'h310a: char_row_bitmap <= 16'b0000001100000000;
		15'h310b: char_row_bitmap <= 16'b0000001110000000;
		15'h310c: char_row_bitmap <= 16'b0000000111000000;
		15'h310d: char_row_bitmap <= 16'b0000000011110000;
		15'h310e: char_row_bitmap <= 16'b0000000000111100;
		15'h310f: char_row_bitmap <= 16'b0000000000111100;
		15'h3110: char_row_bitmap <= 16'b0000000011110000;
		15'h3111: char_row_bitmap <= 16'b0000000111000000;
		15'h3112: char_row_bitmap <= 16'b0000001110000000;
		15'h3113: char_row_bitmap <= 16'b0000001100000000;
		15'h3114: char_row_bitmap <= 16'b0000001100000000;
		15'h3115: char_row_bitmap <= 16'b0000001100000000;
		15'h3116: char_row_bitmap <= 16'b0000001100000000;
		15'h3117: char_row_bitmap <= 16'b0000001100000000;
		15'h3118: char_row_bitmap <= 16'b0000001100000000;
		15'h3119: char_row_bitmap <= 16'b0000001100000000;
		15'h311a: char_row_bitmap <= 16'b0000001100000000;
		15'h311b: char_row_bitmap <= 16'b0000001100000000;
		15'h311c: char_row_bitmap <= 16'b0000001100000000;
		15'h311d: char_row_bitmap <= 16'b0000011100000000;
		15'h311e: char_row_bitmap <= 16'b0000011000000000;
		15'h311f: char_row_bitmap <= 16'b0000111000000000;
		15'h3120: char_row_bitmap <= 16'b0011110000000000;
		15'h3121: char_row_bitmap <= 16'b0011100000000000;
		15'h3122: char_row_bitmap <= 16'b0000000000000000;
		15'h3123: char_row_bitmap <= 16'b0000000000000000;
		15'h3124: char_row_bitmap <= 16'b0000001100000000;
		15'h3125: char_row_bitmap <= 16'b0000001100000000;
		15'h3126: char_row_bitmap <= 16'b0000001100000000;
		15'h3127: char_row_bitmap <= 16'b0000001100000000;
		15'h3128: char_row_bitmap <= 16'b0000001100000000;
		15'h3129: char_row_bitmap <= 16'b0000001100000000;
		15'h312a: char_row_bitmap <= 16'b0000001100000000;
		15'h312b: char_row_bitmap <= 16'b0000001100000000;
		15'h312c: char_row_bitmap <= 16'b0000001100000000;
		15'h312d: char_row_bitmap <= 16'b0000001100000000;
		15'h312e: char_row_bitmap <= 16'b0000001100000000;
		15'h312f: char_row_bitmap <= 16'b0000001100000000;
		15'h3130: char_row_bitmap <= 16'b0000001100000000;
		15'h3131: char_row_bitmap <= 16'b0000001100000000;
		15'h3132: char_row_bitmap <= 16'b0000001100000000;
		15'h3133: char_row_bitmap <= 16'b0000001110000000;
		15'h3134: char_row_bitmap <= 16'b0000000111000000;
		15'h3135: char_row_bitmap <= 16'b0000000011110000;
		15'h3136: char_row_bitmap <= 16'b0000000000111100;
		15'h3137: char_row_bitmap <= 16'b0000000000111100;
		15'h3138: char_row_bitmap <= 16'b0000000011110000;
		15'h3139: char_row_bitmap <= 16'b0000000111000000;
		15'h313a: char_row_bitmap <= 16'b0000001110000000;
		15'h313b: char_row_bitmap <= 16'b0000001100000000;
		15'h313c: char_row_bitmap <= 16'b0000001100000000;
		15'h313d: char_row_bitmap <= 16'b0000001100000000;
		15'h313e: char_row_bitmap <= 16'b0000001100000000;
		15'h313f: char_row_bitmap <= 16'b0000001100000000;
		15'h3140: char_row_bitmap <= 16'b0000001100000000;
		15'h3141: char_row_bitmap <= 16'b0000001100000000;
		15'h3142: char_row_bitmap <= 16'b0000001100000000;
		15'h3143: char_row_bitmap <= 16'b0000001100000000;
		15'h3144: char_row_bitmap <= 16'b0000001100000000;
		15'h3145: char_row_bitmap <= 16'b0000001100000000;
		15'h3146: char_row_bitmap <= 16'b0000001100000000;
		15'h3147: char_row_bitmap <= 16'b0000001100000000;
		15'h3148: char_row_bitmap <= 16'b0000001100000000;
		15'h3149: char_row_bitmap <= 16'b0000001100000000;
		15'h314a: char_row_bitmap <= 16'b0000001100000000;
		15'h314b: char_row_bitmap <= 16'b0000001100000000;
		15'h314c: char_row_bitmap <= 16'b0000000000011100;
		15'h314d: char_row_bitmap <= 16'b0000000000111100;
		15'h314e: char_row_bitmap <= 16'b0000000001110000;
		15'h314f: char_row_bitmap <= 16'b0000000001100000;
		15'h3150: char_row_bitmap <= 16'b0000000011100000;
		15'h3151: char_row_bitmap <= 16'b0000000011000000;
		15'h3152: char_row_bitmap <= 16'b0000000011000000;
		15'h3153: char_row_bitmap <= 16'b0000000011000000;
		15'h3154: char_row_bitmap <= 16'b0000000011000000;
		15'h3155: char_row_bitmap <= 16'b0000000011000000;
		15'h3156: char_row_bitmap <= 16'b0000000011000000;
		15'h3157: char_row_bitmap <= 16'b0000000011000000;
		15'h3158: char_row_bitmap <= 16'b0000000011000000;
		15'h3159: char_row_bitmap <= 16'b0000000011000000;
		15'h315a: char_row_bitmap <= 16'b0000000011000000;
		15'h315b: char_row_bitmap <= 16'b0000000011000000;
		15'h315c: char_row_bitmap <= 16'b0000000011000000;
		15'h315d: char_row_bitmap <= 16'b0000000011000000;
		15'h315e: char_row_bitmap <= 16'b0000000011000000;
		15'h315f: char_row_bitmap <= 16'b0000000011000000;
		15'h3160: char_row_bitmap <= 16'b0000000011000000;
		15'h3161: char_row_bitmap <= 16'b0000000011000000;
		15'h3162: char_row_bitmap <= 16'b0000000011000000;
		15'h3163: char_row_bitmap <= 16'b0000000011000000;
		15'h3164: char_row_bitmap <= 16'b0000000011000000;
		15'h3165: char_row_bitmap <= 16'b0000000011000000;
		15'h3166: char_row_bitmap <= 16'b0000000011000000;
		15'h3167: char_row_bitmap <= 16'b0000000011000000;
		15'h3168: char_row_bitmap <= 16'b0000000011000000;
		15'h3169: char_row_bitmap <= 16'b0000000011000000;
		15'h316a: char_row_bitmap <= 16'b0000000011000000;
		15'h316b: char_row_bitmap <= 16'b0000000011000000;
		15'h316c: char_row_bitmap <= 16'b0000000011000000;
		15'h316d: char_row_bitmap <= 16'b0000000011100000;
		15'h316e: char_row_bitmap <= 16'b0000000001100000;
		15'h316f: char_row_bitmap <= 16'b0000000001110000;
		15'h3170: char_row_bitmap <= 16'b0000000000111100;
		15'h3171: char_row_bitmap <= 16'b0000000000011100;
		15'h3172: char_row_bitmap <= 16'b0000000000000000;
		15'h3173: char_row_bitmap <= 16'b0000000000000000;
		15'h3174: char_row_bitmap <= 16'b0000000011000000;
		15'h3175: char_row_bitmap <= 16'b0000000011000000;
		15'h3176: char_row_bitmap <= 16'b0000000011000000;
		15'h3177: char_row_bitmap <= 16'b0000000011000000;
		15'h3178: char_row_bitmap <= 16'b0000000011000000;
		15'h3179: char_row_bitmap <= 16'b0000000111000000;
		15'h317a: char_row_bitmap <= 16'b0000001110000000;
		15'h317b: char_row_bitmap <= 16'b0000111100000000;
		15'h317c: char_row_bitmap <= 16'b0011110000000000;
		15'h317d: char_row_bitmap <= 16'b0011110000000000;
		15'h317e: char_row_bitmap <= 16'b0000111100000000;
		15'h317f: char_row_bitmap <= 16'b0000001110000000;
		15'h3180: char_row_bitmap <= 16'b0000000111000000;
		15'h3181: char_row_bitmap <= 16'b0000000011000000;
		15'h3182: char_row_bitmap <= 16'b0000000011000000;
		15'h3183: char_row_bitmap <= 16'b0000000011000000;
		15'h3184: char_row_bitmap <= 16'b0000000011000000;
		15'h3185: char_row_bitmap <= 16'b0000000011000000;
		15'h3186: char_row_bitmap <= 16'b0000000011000000;
		15'h3187: char_row_bitmap <= 16'b0000000011000000;
		15'h3188: char_row_bitmap <= 16'b0000000000011100;
		15'h3189: char_row_bitmap <= 16'b0000000000111100;
		15'h318a: char_row_bitmap <= 16'b0000000001110000;
		15'h318b: char_row_bitmap <= 16'b0000000001100000;
		15'h318c: char_row_bitmap <= 16'b0000000011100000;
		15'h318d: char_row_bitmap <= 16'b0000000011000000;
		15'h318e: char_row_bitmap <= 16'b0000000011000000;
		15'h318f: char_row_bitmap <= 16'b0000000011000000;
		15'h3190: char_row_bitmap <= 16'b0000000011000000;
		15'h3191: char_row_bitmap <= 16'b0000000011000000;
		15'h3192: char_row_bitmap <= 16'b0000000011000000;
		15'h3193: char_row_bitmap <= 16'b0000000011000000;
		15'h3194: char_row_bitmap <= 16'b0000000011000000;
		15'h3195: char_row_bitmap <= 16'b0000000011000000;
		15'h3196: char_row_bitmap <= 16'b0000000011000000;
		15'h3197: char_row_bitmap <= 16'b0000000111000000;
		15'h3198: char_row_bitmap <= 16'b0000001110000000;
		15'h3199: char_row_bitmap <= 16'b0000111100000000;
		15'h319a: char_row_bitmap <= 16'b0011110000000000;
		15'h319b: char_row_bitmap <= 16'b0011110000000000;
		15'h319c: char_row_bitmap <= 16'b0000111100000000;
		15'h319d: char_row_bitmap <= 16'b0000001110000000;
		15'h319e: char_row_bitmap <= 16'b0000000111000000;
		15'h319f: char_row_bitmap <= 16'b0000000011000000;
		15'h31a0: char_row_bitmap <= 16'b0000000011000000;
		15'h31a1: char_row_bitmap <= 16'b0000000011000000;
		15'h31a2: char_row_bitmap <= 16'b0000000011000000;
		15'h31a3: char_row_bitmap <= 16'b0000000011000000;
		15'h31a4: char_row_bitmap <= 16'b0000000011000000;
		15'h31a5: char_row_bitmap <= 16'b0000000011000000;
		15'h31a6: char_row_bitmap <= 16'b0000000011000000;
		15'h31a7: char_row_bitmap <= 16'b0000000011000000;
		15'h31a8: char_row_bitmap <= 16'b0000000011000000;
		15'h31a9: char_row_bitmap <= 16'b0000000011100000;
		15'h31aa: char_row_bitmap <= 16'b0000000001100000;
		15'h31ab: char_row_bitmap <= 16'b0000000001110000;
		15'h31ac: char_row_bitmap <= 16'b0000000000111100;
		15'h31ad: char_row_bitmap <= 16'b0000000000011100;
		15'h31ae: char_row_bitmap <= 16'b0000000000000000;
		15'h31af: char_row_bitmap <= 16'b0000000000000000;
		15'h31b0: char_row_bitmap <= 16'b0000000011000000;
		15'h31b1: char_row_bitmap <= 16'b0000000011000000;
		15'h31b2: char_row_bitmap <= 16'b0000000011000000;
		15'h31b3: char_row_bitmap <= 16'b0000000011000000;
		15'h31b4: char_row_bitmap <= 16'b0000000011000000;
		15'h31b5: char_row_bitmap <= 16'b0000000011000000;
		15'h31b6: char_row_bitmap <= 16'b0000000011000000;
		15'h31b7: char_row_bitmap <= 16'b0000000011000000;
		15'h31b8: char_row_bitmap <= 16'b0000000011000000;
		15'h31b9: char_row_bitmap <= 16'b0000000011000000;
		15'h31ba: char_row_bitmap <= 16'b0000000011000000;
		15'h31bb: char_row_bitmap <= 16'b0000000011000000;
		15'h31bc: char_row_bitmap <= 16'b0000000011000000;
		15'h31bd: char_row_bitmap <= 16'b0000000011000000;
		15'h31be: char_row_bitmap <= 16'b0000000011000000;
		15'h31bf: char_row_bitmap <= 16'b0000000111000000;
		15'h31c0: char_row_bitmap <= 16'b0000001110000000;
		15'h31c1: char_row_bitmap <= 16'b0000111100000000;
		15'h31c2: char_row_bitmap <= 16'b0011110000000000;
		15'h31c3: char_row_bitmap <= 16'b0011110000000000;
		15'h31c4: char_row_bitmap <= 16'b0000111100000000;
		15'h31c5: char_row_bitmap <= 16'b0000001110000000;
		15'h31c6: char_row_bitmap <= 16'b0000000111000000;
		15'h31c7: char_row_bitmap <= 16'b0000000011000000;
		15'h31c8: char_row_bitmap <= 16'b0000000011000000;
		15'h31c9: char_row_bitmap <= 16'b0000000011000000;
		15'h31ca: char_row_bitmap <= 16'b0000000011000000;
		15'h31cb: char_row_bitmap <= 16'b0000000011000000;
		15'h31cc: char_row_bitmap <= 16'b0000000011000000;
		15'h31cd: char_row_bitmap <= 16'b0000000011000000;
		15'h31ce: char_row_bitmap <= 16'b0000000011000000;
		15'h31cf: char_row_bitmap <= 16'b0000000011000000;
		15'h31d0: char_row_bitmap <= 16'b0000000011000000;
		15'h31d1: char_row_bitmap <= 16'b0000000011000000;
		15'h31d2: char_row_bitmap <= 16'b0000000011000000;
		15'h31d3: char_row_bitmap <= 16'b0000000011000000;
		15'h31d4: char_row_bitmap <= 16'b0000000011000000;
		15'h31d5: char_row_bitmap <= 16'b0000000011000000;
		15'h31d6: char_row_bitmap <= 16'b0000000011000000;
		15'h31d7: char_row_bitmap <= 16'b0000000011000000;
		15'h31d8: char_row_bitmap <= 16'b0000000011000000;
		15'h31d9: char_row_bitmap <= 16'b0000000011000000;
		15'h31da: char_row_bitmap <= 16'b0000000011000000;
		15'h31db: char_row_bitmap <= 16'b0000000011000000;
		15'h31dc: char_row_bitmap <= 16'b0000000011000000;
		15'h31dd: char_row_bitmap <= 16'b0000000111000000;
		15'h31de: char_row_bitmap <= 16'b0000001110000000;
		15'h31df: char_row_bitmap <= 16'b0000111100000000;
		15'h31e0: char_row_bitmap <= 16'b0011110000000000;
		15'h31e1: char_row_bitmap <= 16'b0011110000000000;
		15'h31e2: char_row_bitmap <= 16'b0000111100000000;
		15'h31e3: char_row_bitmap <= 16'b0000001110000000;
		15'h31e4: char_row_bitmap <= 16'b0000000111000000;
		15'h31e5: char_row_bitmap <= 16'b0000000011100000;
		15'h31e6: char_row_bitmap <= 16'b0000000001100000;
		15'h31e7: char_row_bitmap <= 16'b0000000001110000;
		15'h31e8: char_row_bitmap <= 16'b0000000000111100;
		15'h31e9: char_row_bitmap <= 16'b0000000000011100;
		15'h31ea: char_row_bitmap <= 16'b0000000000000000;
		15'h31eb: char_row_bitmap <= 16'b0000000000000000;
		15'h31ec: char_row_bitmap <= 16'b0000001100000000;
		15'h31ed: char_row_bitmap <= 16'b0000001100000000;
		15'h31ee: char_row_bitmap <= 16'b0000001100000000;
		15'h31ef: char_row_bitmap <= 16'b0000001100000000;
		15'h31f0: char_row_bitmap <= 16'b0000001100000000;
		15'h31f1: char_row_bitmap <= 16'b0000001110000000;
		15'h31f2: char_row_bitmap <= 16'b0000000111000000;
		15'h31f3: char_row_bitmap <= 16'b0000000011110000;
		15'h31f4: char_row_bitmap <= 16'b0000000000111100;
		15'h31f5: char_row_bitmap <= 16'b0000000000111100;
		15'h31f6: char_row_bitmap <= 16'b0000000011110000;
		15'h31f7: char_row_bitmap <= 16'b0000000111000000;
		15'h31f8: char_row_bitmap <= 16'b0000001110000000;
		15'h31f9: char_row_bitmap <= 16'b0000011100000000;
		15'h31fa: char_row_bitmap <= 16'b0000011000000000;
		15'h31fb: char_row_bitmap <= 16'b0000111000000000;
		15'h31fc: char_row_bitmap <= 16'b0011110000000000;
		15'h31fd: char_row_bitmap <= 16'b0011100000000000;
		15'h31fe: char_row_bitmap <= 16'b0000000000000000;
		15'h31ff: char_row_bitmap <= 16'b0000000000000000;
		15'h3200: char_row_bitmap <= 16'b1100000000000000;
		15'h3201: char_row_bitmap <= 16'b1100000000000000;
		15'h3202: char_row_bitmap <= 16'b1100000000000000;
		15'h3203: char_row_bitmap <= 16'b1100000000000000;
		15'h3204: char_row_bitmap <= 16'b1100000000000000;
		15'h3205: char_row_bitmap <= 16'b1100000000000000;
		15'h3206: char_row_bitmap <= 16'b1100000000000000;
		15'h3207: char_row_bitmap <= 16'b1100000000000000;
		15'h3208: char_row_bitmap <= 16'b1100000000000000;
		15'h3209: char_row_bitmap <= 16'b1100000000000000;
		15'h320a: char_row_bitmap <= 16'b1100000000000000;
		15'h320b: char_row_bitmap <= 16'b1100000000000000;
		15'h320c: char_row_bitmap <= 16'b1100000000000000;
		15'h320d: char_row_bitmap <= 16'b1100000000000000;
		15'h320e: char_row_bitmap <= 16'b1100000000000000;
		15'h320f: char_row_bitmap <= 16'b1100000000000000;
		15'h3210: char_row_bitmap <= 16'b1100000000000000;
		15'h3211: char_row_bitmap <= 16'b1100000000000000;
		15'h3212: char_row_bitmap <= 16'b1100000000000000;
		15'h3213: char_row_bitmap <= 16'b1100000000000000;
		15'h3214: char_row_bitmap <= 16'b0011000000000000;
		15'h3215: char_row_bitmap <= 16'b0011000000000000;
		15'h3216: char_row_bitmap <= 16'b0011000000000000;
		15'h3217: char_row_bitmap <= 16'b0011000000000000;
		15'h3218: char_row_bitmap <= 16'b0011000000000000;
		15'h3219: char_row_bitmap <= 16'b0011000000000000;
		15'h321a: char_row_bitmap <= 16'b0011000000000000;
		15'h321b: char_row_bitmap <= 16'b0011000000000000;
		15'h321c: char_row_bitmap <= 16'b0011000000000000;
		15'h321d: char_row_bitmap <= 16'b0011000000000000;
		15'h321e: char_row_bitmap <= 16'b0011000000000000;
		15'h321f: char_row_bitmap <= 16'b0011000000000000;
		15'h3220: char_row_bitmap <= 16'b0011000000000000;
		15'h3221: char_row_bitmap <= 16'b0011000000000000;
		15'h3222: char_row_bitmap <= 16'b0011000000000000;
		15'h3223: char_row_bitmap <= 16'b0011000000000000;
		15'h3224: char_row_bitmap <= 16'b0011000000000000;
		15'h3225: char_row_bitmap <= 16'b0011000000000000;
		15'h3226: char_row_bitmap <= 16'b0011000000000000;
		15'h3227: char_row_bitmap <= 16'b0011000000000000;
		15'h3228: char_row_bitmap <= 16'b0000110000000000;
		15'h3229: char_row_bitmap <= 16'b0000110000000000;
		15'h322a: char_row_bitmap <= 16'b0000110000000000;
		15'h322b: char_row_bitmap <= 16'b0000110000000000;
		15'h322c: char_row_bitmap <= 16'b0000110000000000;
		15'h322d: char_row_bitmap <= 16'b0000110000000000;
		15'h322e: char_row_bitmap <= 16'b0000110000000000;
		15'h322f: char_row_bitmap <= 16'b0000110000000000;
		15'h3230: char_row_bitmap <= 16'b0000110000000000;
		15'h3231: char_row_bitmap <= 16'b0000110000000000;
		15'h3232: char_row_bitmap <= 16'b0000110000000000;
		15'h3233: char_row_bitmap <= 16'b0000110000000000;
		15'h3234: char_row_bitmap <= 16'b0000110000000000;
		15'h3235: char_row_bitmap <= 16'b0000110000000000;
		15'h3236: char_row_bitmap <= 16'b0000110000000000;
		15'h3237: char_row_bitmap <= 16'b0000110000000000;
		15'h3238: char_row_bitmap <= 16'b0000110000000000;
		15'h3239: char_row_bitmap <= 16'b0000110000000000;
		15'h323a: char_row_bitmap <= 16'b0000110000000000;
		15'h323b: char_row_bitmap <= 16'b0000110000000000;
		15'h323c: char_row_bitmap <= 16'b0000001100000000;
		15'h323d: char_row_bitmap <= 16'b0000001100000000;
		15'h323e: char_row_bitmap <= 16'b0000001100000000;
		15'h323f: char_row_bitmap <= 16'b0000001100000000;
		15'h3240: char_row_bitmap <= 16'b0000001100000000;
		15'h3241: char_row_bitmap <= 16'b0000001100000000;
		15'h3242: char_row_bitmap <= 16'b0000001100000000;
		15'h3243: char_row_bitmap <= 16'b0000001100000000;
		15'h3244: char_row_bitmap <= 16'b0000001100000000;
		15'h3245: char_row_bitmap <= 16'b0000001100000000;
		15'h3246: char_row_bitmap <= 16'b0000001100000000;
		15'h3247: char_row_bitmap <= 16'b0000001100000000;
		15'h3248: char_row_bitmap <= 16'b0000001100000000;
		15'h3249: char_row_bitmap <= 16'b0000001100000000;
		15'h324a: char_row_bitmap <= 16'b0000001100000000;
		15'h324b: char_row_bitmap <= 16'b0000001100000000;
		15'h324c: char_row_bitmap <= 16'b0000001100000000;
		15'h324d: char_row_bitmap <= 16'b0000001100000000;
		15'h324e: char_row_bitmap <= 16'b0000001100000000;
		15'h324f: char_row_bitmap <= 16'b0000001100000000;
		15'h3250: char_row_bitmap <= 16'b0000000011000000;
		15'h3251: char_row_bitmap <= 16'b0000000011000000;
		15'h3252: char_row_bitmap <= 16'b0000000011000000;
		15'h3253: char_row_bitmap <= 16'b0000000011000000;
		15'h3254: char_row_bitmap <= 16'b0000000011000000;
		15'h3255: char_row_bitmap <= 16'b0000000011000000;
		15'h3256: char_row_bitmap <= 16'b0000000011000000;
		15'h3257: char_row_bitmap <= 16'b0000000011000000;
		15'h3258: char_row_bitmap <= 16'b0000000011000000;
		15'h3259: char_row_bitmap <= 16'b0000000011000000;
		15'h325a: char_row_bitmap <= 16'b0000000011000000;
		15'h325b: char_row_bitmap <= 16'b0000000011000000;
		15'h325c: char_row_bitmap <= 16'b0000000011000000;
		15'h325d: char_row_bitmap <= 16'b0000000011000000;
		15'h325e: char_row_bitmap <= 16'b0000000011000000;
		15'h325f: char_row_bitmap <= 16'b0000000011000000;
		15'h3260: char_row_bitmap <= 16'b0000000011000000;
		15'h3261: char_row_bitmap <= 16'b0000000011000000;
		15'h3262: char_row_bitmap <= 16'b0000000011000000;
		15'h3263: char_row_bitmap <= 16'b0000000011000000;
		15'h3264: char_row_bitmap <= 16'b0000000000110000;
		15'h3265: char_row_bitmap <= 16'b0000000000110000;
		15'h3266: char_row_bitmap <= 16'b0000000000110000;
		15'h3267: char_row_bitmap <= 16'b0000000000110000;
		15'h3268: char_row_bitmap <= 16'b0000000000110000;
		15'h3269: char_row_bitmap <= 16'b0000000000110000;
		15'h326a: char_row_bitmap <= 16'b0000000000110000;
		15'h326b: char_row_bitmap <= 16'b0000000000110000;
		15'h326c: char_row_bitmap <= 16'b0000000000110000;
		15'h326d: char_row_bitmap <= 16'b0000000000110000;
		15'h326e: char_row_bitmap <= 16'b0000000000110000;
		15'h326f: char_row_bitmap <= 16'b0000000000110000;
		15'h3270: char_row_bitmap <= 16'b0000000000110000;
		15'h3271: char_row_bitmap <= 16'b0000000000110000;
		15'h3272: char_row_bitmap <= 16'b0000000000110000;
		15'h3273: char_row_bitmap <= 16'b0000000000110000;
		15'h3274: char_row_bitmap <= 16'b0000000000110000;
		15'h3275: char_row_bitmap <= 16'b0000000000110000;
		15'h3276: char_row_bitmap <= 16'b0000000000110000;
		15'h3277: char_row_bitmap <= 16'b0000000000110000;
		15'h3278: char_row_bitmap <= 16'b0000000000001100;
		15'h3279: char_row_bitmap <= 16'b0000000000001100;
		15'h327a: char_row_bitmap <= 16'b0000000000001100;
		15'h327b: char_row_bitmap <= 16'b0000000000001100;
		15'h327c: char_row_bitmap <= 16'b0000000000001100;
		15'h327d: char_row_bitmap <= 16'b0000000000001100;
		15'h327e: char_row_bitmap <= 16'b0000000000001100;
		15'h327f: char_row_bitmap <= 16'b0000000000001100;
		15'h3280: char_row_bitmap <= 16'b0000000000001100;
		15'h3281: char_row_bitmap <= 16'b0000000000001100;
		15'h3282: char_row_bitmap <= 16'b0000000000001100;
		15'h3283: char_row_bitmap <= 16'b0000000000001100;
		15'h3284: char_row_bitmap <= 16'b0000000000001100;
		15'h3285: char_row_bitmap <= 16'b0000000000001100;
		15'h3286: char_row_bitmap <= 16'b0000000000001100;
		15'h3287: char_row_bitmap <= 16'b0000000000001100;
		15'h3288: char_row_bitmap <= 16'b0000000000001100;
		15'h3289: char_row_bitmap <= 16'b0000000000001100;
		15'h328a: char_row_bitmap <= 16'b0000000000001100;
		15'h328b: char_row_bitmap <= 16'b0000000000001100;
		15'h328c: char_row_bitmap <= 16'b0000000000000011;
		15'h328d: char_row_bitmap <= 16'b0000000000000011;
		15'h328e: char_row_bitmap <= 16'b0000000000000011;
		15'h328f: char_row_bitmap <= 16'b0000000000000011;
		15'h3290: char_row_bitmap <= 16'b0000000000000011;
		15'h3291: char_row_bitmap <= 16'b0000000000000011;
		15'h3292: char_row_bitmap <= 16'b0000000000000011;
		15'h3293: char_row_bitmap <= 16'b0000000000000011;
		15'h3294: char_row_bitmap <= 16'b0000000000000011;
		15'h3295: char_row_bitmap <= 16'b0000000000000011;
		15'h3296: char_row_bitmap <= 16'b0000000000000011;
		15'h3297: char_row_bitmap <= 16'b0000000000000011;
		15'h3298: char_row_bitmap <= 16'b0000000000000011;
		15'h3299: char_row_bitmap <= 16'b0000000000000011;
		15'h329a: char_row_bitmap <= 16'b0000000000000011;
		15'h329b: char_row_bitmap <= 16'b0000000000000011;
		15'h329c: char_row_bitmap <= 16'b0000000000000011;
		15'h329d: char_row_bitmap <= 16'b0000000000000011;
		15'h329e: char_row_bitmap <= 16'b0000000000000011;
		15'h329f: char_row_bitmap <= 16'b0000000000000011;
		15'h32a0: char_row_bitmap <= 16'b0000000000000011;
		15'h32a1: char_row_bitmap <= 16'b0000000000000011;
		15'h32a2: char_row_bitmap <= 16'b0000000000000011;
		15'h32a3: char_row_bitmap <= 16'b0000000000000011;
		15'h32a4: char_row_bitmap <= 16'b0000000000000111;
		15'h32a5: char_row_bitmap <= 16'b0000000000001111;
		15'h32a6: char_row_bitmap <= 16'b0000000000111110;
		15'h32a7: char_row_bitmap <= 16'b0000000011111100;
		15'h32a8: char_row_bitmap <= 16'b0000001111110000;
		15'h32a9: char_row_bitmap <= 16'b0000111111000000;
		15'h32aa: char_row_bitmap <= 16'b0011111100000000;
		15'h32ab: char_row_bitmap <= 16'b0011111100000000;
		15'h32ac: char_row_bitmap <= 16'b0000111111000000;
		15'h32ad: char_row_bitmap <= 16'b0000001111110000;
		15'h32ae: char_row_bitmap <= 16'b0000000011111100;
		15'h32af: char_row_bitmap <= 16'b0000000000111110;
		15'h32b0: char_row_bitmap <= 16'b0000000000001111;
		15'h32b1: char_row_bitmap <= 16'b0000000000000111;
		15'h32b2: char_row_bitmap <= 16'b0000000000000011;
		15'h32b3: char_row_bitmap <= 16'b0000000000000011;
		15'h32b4: char_row_bitmap <= 16'b1100000000000000;
		15'h32b5: char_row_bitmap <= 16'b1100000000000000;
		15'h32b6: char_row_bitmap <= 16'b1100000000000000;
		15'h32b7: char_row_bitmap <= 16'b1100000000000000;
		15'h32b8: char_row_bitmap <= 16'b1110000000000000;
		15'h32b9: char_row_bitmap <= 16'b1111000000000000;
		15'h32ba: char_row_bitmap <= 16'b0111110000000000;
		15'h32bb: char_row_bitmap <= 16'b0011111100000000;
		15'h32bc: char_row_bitmap <= 16'b0000111111000000;
		15'h32bd: char_row_bitmap <= 16'b0000001111110000;
		15'h32be: char_row_bitmap <= 16'b0000000011111100;
		15'h32bf: char_row_bitmap <= 16'b0000000011111100;
		15'h32c0: char_row_bitmap <= 16'b0000001111110000;
		15'h32c1: char_row_bitmap <= 16'b0000111111000000;
		15'h32c2: char_row_bitmap <= 16'b0011111100000000;
		15'h32c3: char_row_bitmap <= 16'b0111110000000000;
		15'h32c4: char_row_bitmap <= 16'b1111000000000000;
		15'h32c5: char_row_bitmap <= 16'b1110000000000000;
		15'h32c6: char_row_bitmap <= 16'b1100000000000000;
		15'h32c7: char_row_bitmap <= 16'b1100000000000000;
		15'h32c8: char_row_bitmap <= 16'b1100000000001111;
		15'h32c9: char_row_bitmap <= 16'b1110000000011111;
		15'h32ca: char_row_bitmap <= 16'b1111000000111100;
		15'h32cb: char_row_bitmap <= 16'b0111000000111000;
		15'h32cc: char_row_bitmap <= 16'b0011100001110000;
		15'h32cd: char_row_bitmap <= 16'b0011100001110000;
		15'h32ce: char_row_bitmap <= 16'b0001110011100000;
		15'h32cf: char_row_bitmap <= 16'b0001110011100000;
		15'h32d0: char_row_bitmap <= 16'b0000111111000000;
		15'h32d1: char_row_bitmap <= 16'b0000111111000000;
		15'h32d2: char_row_bitmap <= 16'b0000011110000000;
		15'h32d3: char_row_bitmap <= 16'b0000011110000000;
		15'h32d4: char_row_bitmap <= 16'b0000001100000000;
		15'h32d5: char_row_bitmap <= 16'b0000001100000000;
		15'h32d6: char_row_bitmap <= 16'b0000000000000000;
		15'h32d7: char_row_bitmap <= 16'b0000000000000000;
		15'h32d8: char_row_bitmap <= 16'b0000000000000000;
		15'h32d9: char_row_bitmap <= 16'b0000000000000000;
		15'h32da: char_row_bitmap <= 16'b0000000000000000;
		15'h32db: char_row_bitmap <= 16'b0000000000000000;
		15'h32dc: char_row_bitmap <= 16'b0000000000000000;
		15'h32dd: char_row_bitmap <= 16'b0000000000000000;
		15'h32de: char_row_bitmap <= 16'b0000000000000000;
		15'h32df: char_row_bitmap <= 16'b0000000000000000;
		15'h32e0: char_row_bitmap <= 16'b0000000000000000;
		15'h32e1: char_row_bitmap <= 16'b0000000000000000;
		15'h32e2: char_row_bitmap <= 16'b0000001100000000;
		15'h32e3: char_row_bitmap <= 16'b0000001100000000;
		15'h32e4: char_row_bitmap <= 16'b0000011110000000;
		15'h32e5: char_row_bitmap <= 16'b0000011110000000;
		15'h32e6: char_row_bitmap <= 16'b0000111111000000;
		15'h32e7: char_row_bitmap <= 16'b0000111111000000;
		15'h32e8: char_row_bitmap <= 16'b0001110011100000;
		15'h32e9: char_row_bitmap <= 16'b0001110011100000;
		15'h32ea: char_row_bitmap <= 16'b0011100001110000;
		15'h32eb: char_row_bitmap <= 16'b0011100001110000;
		15'h32ec: char_row_bitmap <= 16'b0111000000111000;
		15'h32ed: char_row_bitmap <= 16'b1111000000111100;
		15'h32ee: char_row_bitmap <= 16'b1110000000011111;
		15'h32ef: char_row_bitmap <= 16'b1100000000001111;
		15'h32f0: char_row_bitmap <= 16'b0000000000000011;
		15'h32f1: char_row_bitmap <= 16'b0000000000000011;
		15'h32f2: char_row_bitmap <= 16'b0000000000000011;
		15'h32f3: char_row_bitmap <= 16'b0000000000000011;
		15'h32f4: char_row_bitmap <= 16'b0000000000000011;
		15'h32f5: char_row_bitmap <= 16'b0000000000001111;
		15'h32f6: char_row_bitmap <= 16'b0000000000111111;
		15'h32f7: char_row_bitmap <= 16'b0000000011111111;
		15'h32f8: char_row_bitmap <= 16'b0000001111111111;
		15'h32f9: char_row_bitmap <= 16'b0000111111111111;
		15'h32fa: char_row_bitmap <= 16'b0011111111111111;
		15'h32fb: char_row_bitmap <= 16'b0011111111111111;
		15'h32fc: char_row_bitmap <= 16'b0000111111111111;
		15'h32fd: char_row_bitmap <= 16'b0000001111111111;
		15'h32fe: char_row_bitmap <= 16'b0000000011111111;
		15'h32ff: char_row_bitmap <= 16'b0000000000111111;
		15'h3300: char_row_bitmap <= 16'b0000000000001111;
		15'h3301: char_row_bitmap <= 16'b0000000000000011;
		15'h3302: char_row_bitmap <= 16'b0000000000000011;
		15'h3303: char_row_bitmap <= 16'b0000000000000011;
		15'h3304: char_row_bitmap <= 16'b1100000000000000;
		15'h3305: char_row_bitmap <= 16'b1100000000000000;
		15'h3306: char_row_bitmap <= 16'b1100000000000000;
		15'h3307: char_row_bitmap <= 16'b1100000000000000;
		15'h3308: char_row_bitmap <= 16'b1100000000000000;
		15'h3309: char_row_bitmap <= 16'b1111000000000000;
		15'h330a: char_row_bitmap <= 16'b1111110000000000;
		15'h330b: char_row_bitmap <= 16'b1111111100000000;
		15'h330c: char_row_bitmap <= 16'b1111111111000000;
		15'h330d: char_row_bitmap <= 16'b1111111111110000;
		15'h330e: char_row_bitmap <= 16'b1111111111111100;
		15'h330f: char_row_bitmap <= 16'b1111111111111100;
		15'h3310: char_row_bitmap <= 16'b1111111111110000;
		15'h3311: char_row_bitmap <= 16'b1111111111000000;
		15'h3312: char_row_bitmap <= 16'b1111111100000000;
		15'h3313: char_row_bitmap <= 16'b1111110000000000;
		15'h3314: char_row_bitmap <= 16'b1111000000000000;
		15'h3315: char_row_bitmap <= 16'b1100000000000000;
		15'h3316: char_row_bitmap <= 16'b1100000000000000;
		15'h3317: char_row_bitmap <= 16'b1100000000000000;
		15'h3318: char_row_bitmap <= 16'b1111111111111111;
		15'h3319: char_row_bitmap <= 16'b1111111111111111;
		15'h331a: char_row_bitmap <= 16'b0111111111111000;
		15'h331b: char_row_bitmap <= 16'b0111111111111000;
		15'h331c: char_row_bitmap <= 16'b0011111111110000;
		15'h331d: char_row_bitmap <= 16'b0011111111110000;
		15'h331e: char_row_bitmap <= 16'b0001111111100000;
		15'h331f: char_row_bitmap <= 16'b0001111111100000;
		15'h3320: char_row_bitmap <= 16'b0000111111000000;
		15'h3321: char_row_bitmap <= 16'b0000111111000000;
		15'h3322: char_row_bitmap <= 16'b0000011110000000;
		15'h3323: char_row_bitmap <= 16'b0000011110000000;
		15'h3324: char_row_bitmap <= 16'b0000001100000000;
		15'h3325: char_row_bitmap <= 16'b0000001100000000;
		15'h3326: char_row_bitmap <= 16'b0000000000000000;
		15'h3327: char_row_bitmap <= 16'b0000000000000000;
		15'h3328: char_row_bitmap <= 16'b0000000000000000;
		15'h3329: char_row_bitmap <= 16'b0000000000000000;
		15'h332a: char_row_bitmap <= 16'b0000000000000000;
		15'h332b: char_row_bitmap <= 16'b0000000000000000;
		15'h332c: char_row_bitmap <= 16'b0000000000000000;
		15'h332d: char_row_bitmap <= 16'b0000000000000000;
		15'h332e: char_row_bitmap <= 16'b0000000000000000;
		15'h332f: char_row_bitmap <= 16'b0000000000000000;
		15'h3330: char_row_bitmap <= 16'b0000000000000000;
		15'h3331: char_row_bitmap <= 16'b0000000000000000;
		15'h3332: char_row_bitmap <= 16'b0000001100000000;
		15'h3333: char_row_bitmap <= 16'b0000001100000000;
		15'h3334: char_row_bitmap <= 16'b0000011110000000;
		15'h3335: char_row_bitmap <= 16'b0000011110000000;
		15'h3336: char_row_bitmap <= 16'b0000111111000000;
		15'h3337: char_row_bitmap <= 16'b0000111111000000;
		15'h3338: char_row_bitmap <= 16'b0001111111100000;
		15'h3339: char_row_bitmap <= 16'b0001111111100000;
		15'h333a: char_row_bitmap <= 16'b0011111111110000;
		15'h333b: char_row_bitmap <= 16'b0011111111110000;
		15'h333c: char_row_bitmap <= 16'b0111111111111000;
		15'h333d: char_row_bitmap <= 16'b0111111111111000;
		15'h333e: char_row_bitmap <= 16'b1111111111111111;
		15'h333f: char_row_bitmap <= 16'b1111111111111111;
		15'h3340: char_row_bitmap <= 16'b1111111111111111;
		15'h3341: char_row_bitmap <= 16'b1111111111111111;
		15'h3342: char_row_bitmap <= 16'b0000000000000000;
		15'h3343: char_row_bitmap <= 16'b0000000000000000;
		15'h3344: char_row_bitmap <= 16'b0000000000000000;
		15'h3345: char_row_bitmap <= 16'b0000000000000000;
		15'h3346: char_row_bitmap <= 16'b0000000000000000;
		15'h3347: char_row_bitmap <= 16'b0000000000000000;
		15'h3348: char_row_bitmap <= 16'b0000000000000000;
		15'h3349: char_row_bitmap <= 16'b0000000000000000;
		15'h334a: char_row_bitmap <= 16'b0000000000000000;
		15'h334b: char_row_bitmap <= 16'b0000000000000000;
		15'h334c: char_row_bitmap <= 16'b0000000000000000;
		15'h334d: char_row_bitmap <= 16'b0000000000000000;
		15'h334e: char_row_bitmap <= 16'b0000000000000000;
		15'h334f: char_row_bitmap <= 16'b0000000000000000;
		15'h3350: char_row_bitmap <= 16'b0000000000000000;
		15'h3351: char_row_bitmap <= 16'b0000000000000000;
		15'h3352: char_row_bitmap <= 16'b0000000000000000;
		15'h3353: char_row_bitmap <= 16'b0000000000000000;
		15'h3354: char_row_bitmap <= 16'b0000000000000000;
		15'h3355: char_row_bitmap <= 16'b0000000000000000;
		15'h3356: char_row_bitmap <= 16'b1111111111111111;
		15'h3357: char_row_bitmap <= 16'b1111111111111111;
		15'h3358: char_row_bitmap <= 16'b0000000000000000;
		15'h3359: char_row_bitmap <= 16'b0000000000000000;
		15'h335a: char_row_bitmap <= 16'b0000000000000000;
		15'h335b: char_row_bitmap <= 16'b0000000000000000;
		15'h335c: char_row_bitmap <= 16'b0000000000000000;
		15'h335d: char_row_bitmap <= 16'b0000000000000000;
		15'h335e: char_row_bitmap <= 16'b0000000000000000;
		15'h335f: char_row_bitmap <= 16'b0000000000000000;
		15'h3360: char_row_bitmap <= 16'b0000000000000000;
		15'h3361: char_row_bitmap <= 16'b0000000000000000;
		15'h3362: char_row_bitmap <= 16'b0000000000000000;
		15'h3363: char_row_bitmap <= 16'b0000000000000000;
		15'h3364: char_row_bitmap <= 16'b0000000000000000;
		15'h3365: char_row_bitmap <= 16'b0000000000000000;
		15'h3366: char_row_bitmap <= 16'b0000000000000000;
		15'h3367: char_row_bitmap <= 16'b0000000000000000;
		15'h3368: char_row_bitmap <= 16'b0000000000000000;
		15'h3369: char_row_bitmap <= 16'b0000000000000000;
		15'h336a: char_row_bitmap <= 16'b0000000000000000;
		15'h336b: char_row_bitmap <= 16'b0000000000000000;
		15'h336c: char_row_bitmap <= 16'b1111111111111111;
		15'h336d: char_row_bitmap <= 16'b1111111111111111;
		15'h336e: char_row_bitmap <= 16'b0000000000000000;
		15'h336f: char_row_bitmap <= 16'b0000000000000000;
		15'h3370: char_row_bitmap <= 16'b0000000000000000;
		15'h3371: char_row_bitmap <= 16'b0000000000000000;
		15'h3372: char_row_bitmap <= 16'b0000000000000000;
		15'h3373: char_row_bitmap <= 16'b0000000000000000;
		15'h3374: char_row_bitmap <= 16'b0000000000000000;
		15'h3375: char_row_bitmap <= 16'b0000000000000000;
		15'h3376: char_row_bitmap <= 16'b0000000000000000;
		15'h3377: char_row_bitmap <= 16'b0000000000000000;
		15'h3378: char_row_bitmap <= 16'b0000000000000000;
		15'h3379: char_row_bitmap <= 16'b0000000000000000;
		15'h337a: char_row_bitmap <= 16'b0000000000000000;
		15'h337b: char_row_bitmap <= 16'b0000000000000000;
		15'h337c: char_row_bitmap <= 16'b0000000000000000;
		15'h337d: char_row_bitmap <= 16'b0000000000000000;
		15'h337e: char_row_bitmap <= 16'b0000000000000000;
		15'h337f: char_row_bitmap <= 16'b0000000000000000;
		15'h3380: char_row_bitmap <= 16'b0000000000000000;
		15'h3381: char_row_bitmap <= 16'b0000000000000000;
		15'h3382: char_row_bitmap <= 16'b1111111111111111;
		15'h3383: char_row_bitmap <= 16'b1111111111111111;
		15'h3384: char_row_bitmap <= 16'b0000000000000000;
		15'h3385: char_row_bitmap <= 16'b0000000000000000;
		15'h3386: char_row_bitmap <= 16'b0000000000000000;
		15'h3387: char_row_bitmap <= 16'b0000000000000000;
		15'h3388: char_row_bitmap <= 16'b0000000000000000;
		15'h3389: char_row_bitmap <= 16'b0000000000000000;
		15'h338a: char_row_bitmap <= 16'b0000000000000000;
		15'h338b: char_row_bitmap <= 16'b0000000000000000;
		15'h338c: char_row_bitmap <= 16'b0000000000000000;
		15'h338d: char_row_bitmap <= 16'b0000000000000000;
		15'h338e: char_row_bitmap <= 16'b0000000000000000;
		15'h338f: char_row_bitmap <= 16'b0000000000000000;
		15'h3390: char_row_bitmap <= 16'b0000000000000000;
		15'h3391: char_row_bitmap <= 16'b0000000000000000;
		15'h3392: char_row_bitmap <= 16'b0000000000000000;
		15'h3393: char_row_bitmap <= 16'b0000000000000000;
		15'h3394: char_row_bitmap <= 16'b0000000000000000;
		15'h3395: char_row_bitmap <= 16'b0000000000000000;
		15'h3396: char_row_bitmap <= 16'b0000000000000000;
		15'h3397: char_row_bitmap <= 16'b0000000000000000;
		15'h3398: char_row_bitmap <= 16'b1111111111111111;
		15'h3399: char_row_bitmap <= 16'b1111111111111111;
		15'h339a: char_row_bitmap <= 16'b0000000000000000;
		15'h339b: char_row_bitmap <= 16'b0000000000000000;
		15'h339c: char_row_bitmap <= 16'b0000000000000000;
		15'h339d: char_row_bitmap <= 16'b0000000000000000;
		15'h339e: char_row_bitmap <= 16'b0000000000000000;
		15'h339f: char_row_bitmap <= 16'b0000000000000000;
		15'h33a0: char_row_bitmap <= 16'b0000000000000000;
		15'h33a1: char_row_bitmap <= 16'b0000000000000000;
		15'h33a2: char_row_bitmap <= 16'b0000000000000000;
		15'h33a3: char_row_bitmap <= 16'b0000000000000000;
		15'h33a4: char_row_bitmap <= 16'b0000000000000000;
		15'h33a5: char_row_bitmap <= 16'b0000000000000000;
		15'h33a6: char_row_bitmap <= 16'b0000000000000000;
		15'h33a7: char_row_bitmap <= 16'b0000000000000000;
		15'h33a8: char_row_bitmap <= 16'b0000000000000000;
		15'h33a9: char_row_bitmap <= 16'b0000000000000000;
		15'h33aa: char_row_bitmap <= 16'b0000000000000000;
		15'h33ab: char_row_bitmap <= 16'b0000000000000000;
		15'h33ac: char_row_bitmap <= 16'b0000000000000000;
		15'h33ad: char_row_bitmap <= 16'b0000000000000000;
		15'h33ae: char_row_bitmap <= 16'b1111111111111111;
		15'h33af: char_row_bitmap <= 16'b1111111111111111;
		15'h33b0: char_row_bitmap <= 16'b0000000000000000;
		15'h33b1: char_row_bitmap <= 16'b0000000000000000;
		15'h33b2: char_row_bitmap <= 16'b0000000000000000;
		15'h33b3: char_row_bitmap <= 16'b0000000000000000;
		15'h33b4: char_row_bitmap <= 16'b0000000000000000;
		15'h33b5: char_row_bitmap <= 16'b0000000000000000;
		15'h33b6: char_row_bitmap <= 16'b0000000000000000;
		15'h33b7: char_row_bitmap <= 16'b0000000000000000;
		15'h33b8: char_row_bitmap <= 16'b0000000000000000;
		15'h33b9: char_row_bitmap <= 16'b0000000000000000;
		15'h33ba: char_row_bitmap <= 16'b0000000000000000;
		15'h33bb: char_row_bitmap <= 16'b0000000000000000;
		15'h33bc: char_row_bitmap <= 16'b0000000000000000;
		15'h33bd: char_row_bitmap <= 16'b0000000000000000;
		15'h33be: char_row_bitmap <= 16'b0000000000000000;
		15'h33bf: char_row_bitmap <= 16'b0000000000000000;
		15'h33c0: char_row_bitmap <= 16'b0000000000000000;
		15'h33c1: char_row_bitmap <= 16'b0000000000000000;
		15'h33c2: char_row_bitmap <= 16'b0000000000000000;
		15'h33c3: char_row_bitmap <= 16'b0000000000000000;
		15'h33c4: char_row_bitmap <= 16'b1111111111111111;
		15'h33c5: char_row_bitmap <= 16'b1111111111111111;
		15'h33c6: char_row_bitmap <= 16'b0000000000000000;
		15'h33c7: char_row_bitmap <= 16'b0000000000000000;
		15'h33c8: char_row_bitmap <= 16'b0000000000000000;
		15'h33c9: char_row_bitmap <= 16'b0000000000000000;
		15'h33ca: char_row_bitmap <= 16'b0000000000000000;
		15'h33cb: char_row_bitmap <= 16'b0000000000000000;
		15'h33cc: char_row_bitmap <= 16'b0000000000000000;
		15'h33cd: char_row_bitmap <= 16'b0000000000000000;
		15'h33ce: char_row_bitmap <= 16'b0000000000000000;
		15'h33cf: char_row_bitmap <= 16'b0000000000000000;
		15'h33d0: char_row_bitmap <= 16'b0000000000000000;
		15'h33d1: char_row_bitmap <= 16'b0000000000000000;
		15'h33d2: char_row_bitmap <= 16'b0000000000000000;
		15'h33d3: char_row_bitmap <= 16'b0000000000000000;
		15'h33d4: char_row_bitmap <= 16'b0000000000000000;
		15'h33d5: char_row_bitmap <= 16'b0000000000000000;
		15'h33d6: char_row_bitmap <= 16'b0000000000000000;
		15'h33d7: char_row_bitmap <= 16'b0000000000000000;
		15'h33d8: char_row_bitmap <= 16'b0000000000000000;
		15'h33d9: char_row_bitmap <= 16'b0000000000000000;
		15'h33da: char_row_bitmap <= 16'b1111111111111111;
		15'h33db: char_row_bitmap <= 16'b1111111111111111;
		15'h33dc: char_row_bitmap <= 16'b0000000000000000;
		15'h33dd: char_row_bitmap <= 16'b0000000000000000;
		15'h33de: char_row_bitmap <= 16'b0000000000000000;
		15'h33df: char_row_bitmap <= 16'b0000000000000000;
		15'h33e0: char_row_bitmap <= 16'b0000000000000000;
		15'h33e1: char_row_bitmap <= 16'b0000000000000000;
		15'h33e2: char_row_bitmap <= 16'b0000000000000000;
		15'h33e3: char_row_bitmap <= 16'b0000000000000000;
		15'h33e4: char_row_bitmap <= 16'b0000000000000000;
		15'h33e5: char_row_bitmap <= 16'b0000000000000000;
		15'h33e6: char_row_bitmap <= 16'b0000000000000000;
		15'h33e7: char_row_bitmap <= 16'b0000000000000000;
		15'h33e8: char_row_bitmap <= 16'b0000000000000000;
		15'h33e9: char_row_bitmap <= 16'b0000000000000000;
		15'h33ea: char_row_bitmap <= 16'b0000000000000000;
		15'h33eb: char_row_bitmap <= 16'b0000000000000000;
		15'h33ec: char_row_bitmap <= 16'b0000000000000000;
		15'h33ed: char_row_bitmap <= 16'b0000000000000000;
		15'h33ee: char_row_bitmap <= 16'b0000000000000000;
		15'h33ef: char_row_bitmap <= 16'b0000000000000000;
		15'h33f0: char_row_bitmap <= 16'b1111111111111111;
		15'h33f1: char_row_bitmap <= 16'b1111111111111111;
		15'h33f2: char_row_bitmap <= 16'b0000000000000000;
		15'h33f3: char_row_bitmap <= 16'b0000000000000000;
		15'h33f4: char_row_bitmap <= 16'b0000000000000000;
		15'h33f5: char_row_bitmap <= 16'b0000000000000000;
		15'h33f6: char_row_bitmap <= 16'b0000000000000000;
		15'h33f7: char_row_bitmap <= 16'b0000000000000000;
		15'h33f8: char_row_bitmap <= 16'b0000000000000000;
		15'h33f9: char_row_bitmap <= 16'b0000000000000000;
		15'h33fa: char_row_bitmap <= 16'b0000000000000000;
		15'h33fb: char_row_bitmap <= 16'b0000000000000000;
		15'h33fc: char_row_bitmap <= 16'b0000000000000000;
		15'h33fd: char_row_bitmap <= 16'b0000000000000000;
		15'h33fe: char_row_bitmap <= 16'b0000000000000000;
		15'h33ff: char_row_bitmap <= 16'b0000000000000000;
		15'h3400: char_row_bitmap <= 16'b0000000000000000;
		15'h3401: char_row_bitmap <= 16'b0000000000000000;
		15'h3402: char_row_bitmap <= 16'b0000000000000000;
		15'h3403: char_row_bitmap <= 16'b0000000000000000;
		15'h3404: char_row_bitmap <= 16'b0000000000000000;
		15'h3405: char_row_bitmap <= 16'b0000000000000000;
		15'h3406: char_row_bitmap <= 16'b1111111111111111;
		15'h3407: char_row_bitmap <= 16'b1111111111111111;
		15'h3408: char_row_bitmap <= 16'b0000000000000000;
		15'h3409: char_row_bitmap <= 16'b0000000000000000;
		15'h340a: char_row_bitmap <= 16'b0000000000000000;
		15'h340b: char_row_bitmap <= 16'b0000000000000000;
		15'h340c: char_row_bitmap <= 16'b0000000000000000;
		15'h340d: char_row_bitmap <= 16'b0000000000000000;
		15'h340e: char_row_bitmap <= 16'b0000000000000000;
		15'h340f: char_row_bitmap <= 16'b0000000000000000;
		15'h3410: char_row_bitmap <= 16'b0000000000000000;
		15'h3411: char_row_bitmap <= 16'b0000000000000000;
		15'h3412: char_row_bitmap <= 16'b0000000000000000;
		15'h3413: char_row_bitmap <= 16'b0000000110000000;
		15'h3414: char_row_bitmap <= 16'b0000001111000000;
		15'h3415: char_row_bitmap <= 16'b0000011111100000;
		15'h3416: char_row_bitmap <= 16'b0000111111110000;
		15'h3417: char_row_bitmap <= 16'b0001111111111000;
		15'h3418: char_row_bitmap <= 16'b0011111111111100;
		15'h3419: char_row_bitmap <= 16'b0011111111111100;
		15'h341a: char_row_bitmap <= 16'b0000001111000000;
		15'h341b: char_row_bitmap <= 16'b0000001111000000;
		15'h341c: char_row_bitmap <= 16'b0000000000000000;
		15'h341d: char_row_bitmap <= 16'b0000000000000000;
		15'h341e: char_row_bitmap <= 16'b0000000000000000;
		15'h341f: char_row_bitmap <= 16'b0000000000000000;
		15'h3420: char_row_bitmap <= 16'b0011000000000000;
		15'h3421: char_row_bitmap <= 16'b0011100000000000;
		15'h3422: char_row_bitmap <= 16'b0011110000000000;
		15'h3423: char_row_bitmap <= 16'b0011111000000000;
		15'h3424: char_row_bitmap <= 16'b1111111100000000;
		15'h3425: char_row_bitmap <= 16'b1111111110000000;
		15'h3426: char_row_bitmap <= 16'b1111111110000000;
		15'h3427: char_row_bitmap <= 16'b1111111100000000;
		15'h3428: char_row_bitmap <= 16'b0011111000000000;
		15'h3429: char_row_bitmap <= 16'b0011110000000000;
		15'h342a: char_row_bitmap <= 16'b0011100000000000;
		15'h342b: char_row_bitmap <= 16'b0011000000000000;
		15'h342c: char_row_bitmap <= 16'b0000000000000000;
		15'h342d: char_row_bitmap <= 16'b0000000000000000;
		15'h342e: char_row_bitmap <= 16'b0000000000000000;
		15'h342f: char_row_bitmap <= 16'b0000000000000000;
		15'h3430: char_row_bitmap <= 16'b0000001111000000;
		15'h3431: char_row_bitmap <= 16'b0000001111000000;
		15'h3432: char_row_bitmap <= 16'b0011111111111100;
		15'h3433: char_row_bitmap <= 16'b0011111111111100;
		15'h3434: char_row_bitmap <= 16'b0001111111111000;
		15'h3435: char_row_bitmap <= 16'b0000111111110000;
		15'h3436: char_row_bitmap <= 16'b0000011111100000;
		15'h3437: char_row_bitmap <= 16'b0000001111000000;
		15'h3438: char_row_bitmap <= 16'b0000000110000000;
		15'h3439: char_row_bitmap <= 16'b0000000000000000;
		15'h343a: char_row_bitmap <= 16'b0000000000000000;
		15'h343b: char_row_bitmap <= 16'b0000000000000000;
		15'h343c: char_row_bitmap <= 16'b0000000000000000;
		15'h343d: char_row_bitmap <= 16'b0000000000000000;
		15'h343e: char_row_bitmap <= 16'b0000000000000000;
		15'h343f: char_row_bitmap <= 16'b0000000000000000;
		15'h3440: char_row_bitmap <= 16'b0000000000000000;
		15'h3441: char_row_bitmap <= 16'b0000000000000000;
		15'h3442: char_row_bitmap <= 16'b0000000000000000;
		15'h3443: char_row_bitmap <= 16'b0000000000000000;
		15'h3444: char_row_bitmap <= 16'b0000000000000000;
		15'h3445: char_row_bitmap <= 16'b0000000000000000;
		15'h3446: char_row_bitmap <= 16'b0000000000000000;
		15'h3447: char_row_bitmap <= 16'b0000000000000000;
		15'h3448: char_row_bitmap <= 16'b0000000000001100;
		15'h3449: char_row_bitmap <= 16'b0000000000011100;
		15'h344a: char_row_bitmap <= 16'b0000000000111100;
		15'h344b: char_row_bitmap <= 16'b0000000001111100;
		15'h344c: char_row_bitmap <= 16'b0000000011111111;
		15'h344d: char_row_bitmap <= 16'b0000000111111111;
		15'h344e: char_row_bitmap <= 16'b0000000111111111;
		15'h344f: char_row_bitmap <= 16'b0000000011111111;
		15'h3450: char_row_bitmap <= 16'b0000000001111100;
		15'h3451: char_row_bitmap <= 16'b0000000000111100;
		15'h3452: char_row_bitmap <= 16'b0000000000011100;
		15'h3453: char_row_bitmap <= 16'b0000000000001100;
		15'h3454: char_row_bitmap <= 16'b0000000000000000;
		15'h3455: char_row_bitmap <= 16'b0000000000000000;
		15'h3456: char_row_bitmap <= 16'b0000000000000000;
		15'h3457: char_row_bitmap <= 16'b0000000000000000;
		15'h3458: char_row_bitmap <= 16'b0000000000000000;
		15'h3459: char_row_bitmap <= 16'b0000000000000000;
		15'h345a: char_row_bitmap <= 16'b0000000000000000;
		15'h345b: char_row_bitmap <= 16'b0000000000000000;
		15'h345c: char_row_bitmap <= 16'b0000011001100000;
		15'h345d: char_row_bitmap <= 16'b0000111001110000;
		15'h345e: char_row_bitmap <= 16'b0001111001111000;
		15'h345f: char_row_bitmap <= 16'b0011111001111100;
		15'h3460: char_row_bitmap <= 16'b0111111111111110;
		15'h3461: char_row_bitmap <= 16'b1111111111111111;
		15'h3462: char_row_bitmap <= 16'b1111111111111111;
		15'h3463: char_row_bitmap <= 16'b0111111111111110;
		15'h3464: char_row_bitmap <= 16'b0011111001111100;
		15'h3465: char_row_bitmap <= 16'b0001111001111000;
		15'h3466: char_row_bitmap <= 16'b0000111001110000;
		15'h3467: char_row_bitmap <= 16'b0000011001100000;
		15'h3468: char_row_bitmap <= 16'b0000000000000000;
		15'h3469: char_row_bitmap <= 16'b0000000000000000;
		15'h346a: char_row_bitmap <= 16'b0000000000000000;
		15'h346b: char_row_bitmap <= 16'b0000000000000000;
		15'h346c: char_row_bitmap <= 16'b0000000000000000;
		15'h346d: char_row_bitmap <= 16'b0000000110000000;
		15'h346e: char_row_bitmap <= 16'b0000001111000000;
		15'h346f: char_row_bitmap <= 16'b0000011111100000;
		15'h3470: char_row_bitmap <= 16'b0000111111110000;
		15'h3471: char_row_bitmap <= 16'b0001111111111000;
		15'h3472: char_row_bitmap <= 16'b0011111111111100;
		15'h3473: char_row_bitmap <= 16'b0011111111111100;
		15'h3474: char_row_bitmap <= 16'b0000001111000000;
		15'h3475: char_row_bitmap <= 16'b0000001111000000;
		15'h3476: char_row_bitmap <= 16'b0000001111000000;
		15'h3477: char_row_bitmap <= 16'b0000001111000000;
		15'h3478: char_row_bitmap <= 16'b0011111111111100;
		15'h3479: char_row_bitmap <= 16'b0011111111111100;
		15'h347a: char_row_bitmap <= 16'b0001111111111000;
		15'h347b: char_row_bitmap <= 16'b0000111111110000;
		15'h347c: char_row_bitmap <= 16'b0000011111100000;
		15'h347d: char_row_bitmap <= 16'b0000001111000000;
		15'h347e: char_row_bitmap <= 16'b0000000110000000;
		15'h347f: char_row_bitmap <= 16'b0000000000000000;
		15'h3480: char_row_bitmap <= 16'b0000000000000000;
		15'h3481: char_row_bitmap <= 16'b0000000000000000;
		15'h3482: char_row_bitmap <= 16'b0000000000000000;
		15'h3483: char_row_bitmap <= 16'b0000000000000000;
		15'h3484: char_row_bitmap <= 16'b0000000000000000;
		15'h3485: char_row_bitmap <= 16'b0000000000000000;
		15'h3486: char_row_bitmap <= 16'b0000000000000000;
		15'h3487: char_row_bitmap <= 16'b0000000000000000;
		15'h3488: char_row_bitmap <= 16'b0000000000000000;
		15'h3489: char_row_bitmap <= 16'b0000000000000000;
		15'h348a: char_row_bitmap <= 16'b0000000000000000;
		15'h348b: char_row_bitmap <= 16'b0000000000000000;
		15'h348c: char_row_bitmap <= 16'b0000000000000000;
		15'h348d: char_row_bitmap <= 16'b0000000000000000;
		15'h348e: char_row_bitmap <= 16'b1000000000000000;
		15'h348f: char_row_bitmap <= 16'b1100000000000000;
		15'h3490: char_row_bitmap <= 16'b1110000000000000;
		15'h3491: char_row_bitmap <= 16'b1111100000000000;
		15'h3492: char_row_bitmap <= 16'b1111110000000000;
		15'h3493: char_row_bitmap <= 16'b1111111100000000;
		15'h3494: char_row_bitmap <= 16'b0000000000000000;
		15'h3495: char_row_bitmap <= 16'b0000000000000000;
		15'h3496: char_row_bitmap <= 16'b0000000000000000;
		15'h3497: char_row_bitmap <= 16'b0000000000000000;
		15'h3498: char_row_bitmap <= 16'b0000000000000000;
		15'h3499: char_row_bitmap <= 16'b0000000000000000;
		15'h349a: char_row_bitmap <= 16'b0000000000000000;
		15'h349b: char_row_bitmap <= 16'b0000000000000000;
		15'h349c: char_row_bitmap <= 16'b0000000000000000;
		15'h349d: char_row_bitmap <= 16'b0000000000000000;
		15'h349e: char_row_bitmap <= 16'b0000000000000000;
		15'h349f: char_row_bitmap <= 16'b0000000000000000;
		15'h34a0: char_row_bitmap <= 16'b0000000000000000;
		15'h34a1: char_row_bitmap <= 16'b0000000000000000;
		15'h34a2: char_row_bitmap <= 16'b1100000000000000;
		15'h34a3: char_row_bitmap <= 16'b1111000000000000;
		15'h34a4: char_row_bitmap <= 16'b1111111000000000;
		15'h34a5: char_row_bitmap <= 16'b1111111111000000;
		15'h34a6: char_row_bitmap <= 16'b1111111111111000;
		15'h34a7: char_row_bitmap <= 16'b1111111111111110;
		15'h34a8: char_row_bitmap <= 16'b0000000000000000;
		15'h34a9: char_row_bitmap <= 16'b0000000000000000;
		15'h34aa: char_row_bitmap <= 16'b0000000000000000;
		15'h34ab: char_row_bitmap <= 16'b0000000000000000;
		15'h34ac: char_row_bitmap <= 16'b0000000000000000;
		15'h34ad: char_row_bitmap <= 16'b0000000000000000;
		15'h34ae: char_row_bitmap <= 16'b1000000000000000;
		15'h34af: char_row_bitmap <= 16'b1000000000000000;
		15'h34b0: char_row_bitmap <= 16'b1100000000000000;
		15'h34b1: char_row_bitmap <= 16'b1100000000000000;
		15'h34b2: char_row_bitmap <= 16'b1110000000000000;
		15'h34b3: char_row_bitmap <= 16'b1110000000000000;
		15'h34b4: char_row_bitmap <= 16'b1111000000000000;
		15'h34b5: char_row_bitmap <= 16'b1111000000000000;
		15'h34b6: char_row_bitmap <= 16'b1111100000000000;
		15'h34b7: char_row_bitmap <= 16'b1111100000000000;
		15'h34b8: char_row_bitmap <= 16'b1111110000000000;
		15'h34b9: char_row_bitmap <= 16'b1111111000000000;
		15'h34ba: char_row_bitmap <= 16'b1111111000000000;
		15'h34bb: char_row_bitmap <= 16'b1111111100000000;
		15'h34bc: char_row_bitmap <= 16'b0000000000000000;
		15'h34bd: char_row_bitmap <= 16'b0000000000000000;
		15'h34be: char_row_bitmap <= 16'b0000000000000000;
		15'h34bf: char_row_bitmap <= 16'b0000000000000000;
		15'h34c0: char_row_bitmap <= 16'b0000000000000000;
		15'h34c1: char_row_bitmap <= 16'b0000000000000000;
		15'h34c2: char_row_bitmap <= 16'b0000000000000000;
		15'h34c3: char_row_bitmap <= 16'b1000000000000000;
		15'h34c4: char_row_bitmap <= 16'b1100000000000000;
		15'h34c5: char_row_bitmap <= 16'b1111000000000000;
		15'h34c6: char_row_bitmap <= 16'b1111100000000000;
		15'h34c7: char_row_bitmap <= 16'b1111110000000000;
		15'h34c8: char_row_bitmap <= 16'b1111111000000000;
		15'h34c9: char_row_bitmap <= 16'b1111111110000000;
		15'h34ca: char_row_bitmap <= 16'b1111111111000000;
		15'h34cb: char_row_bitmap <= 16'b1111111111100000;
		15'h34cc: char_row_bitmap <= 16'b1111111111110000;
		15'h34cd: char_row_bitmap <= 16'b1111111111111000;
		15'h34ce: char_row_bitmap <= 16'b1111111111111100;
		15'h34cf: char_row_bitmap <= 16'b1111111111111111;
		15'h34d0: char_row_bitmap <= 16'b1000000000000000;
		15'h34d1: char_row_bitmap <= 16'b1000000000000000;
		15'h34d2: char_row_bitmap <= 16'b1100000000000000;
		15'h34d3: char_row_bitmap <= 16'b1100000000000000;
		15'h34d4: char_row_bitmap <= 16'b1100000000000000;
		15'h34d5: char_row_bitmap <= 16'b1110000000000000;
		15'h34d6: char_row_bitmap <= 16'b1110000000000000;
		15'h34d7: char_row_bitmap <= 16'b1110000000000000;
		15'h34d8: char_row_bitmap <= 16'b1111000000000000;
		15'h34d9: char_row_bitmap <= 16'b1111000000000000;
		15'h34da: char_row_bitmap <= 16'b1111000000000000;
		15'h34db: char_row_bitmap <= 16'b1111100000000000;
		15'h34dc: char_row_bitmap <= 16'b1111100000000000;
		15'h34dd: char_row_bitmap <= 16'b1111100000000000;
		15'h34de: char_row_bitmap <= 16'b1111110000000000;
		15'h34df: char_row_bitmap <= 16'b1111110000000000;
		15'h34e0: char_row_bitmap <= 16'b1111111000000000;
		15'h34e1: char_row_bitmap <= 16'b1111111000000000;
		15'h34e2: char_row_bitmap <= 16'b1111111000000000;
		15'h34e3: char_row_bitmap <= 16'b1111111100000000;
		15'h34e4: char_row_bitmap <= 16'b1000000000000000;
		15'h34e5: char_row_bitmap <= 16'b1100000000000000;
		15'h34e6: char_row_bitmap <= 16'b1100000000000000;
		15'h34e7: char_row_bitmap <= 16'b1110000000000000;
		15'h34e8: char_row_bitmap <= 16'b1111000000000000;
		15'h34e9: char_row_bitmap <= 16'b1111000000000000;
		15'h34ea: char_row_bitmap <= 16'b1111100000000000;
		15'h34eb: char_row_bitmap <= 16'b1111110000000000;
		15'h34ec: char_row_bitmap <= 16'b1111111000000000;
		15'h34ed: char_row_bitmap <= 16'b1111111100000000;
		15'h34ee: char_row_bitmap <= 16'b1111111100000000;
		15'h34ef: char_row_bitmap <= 16'b1111111110000000;
		15'h34f0: char_row_bitmap <= 16'b1111111111000000;
		15'h34f1: char_row_bitmap <= 16'b1111111111100000;
		15'h34f2: char_row_bitmap <= 16'b1111111111110000;
		15'h34f3: char_row_bitmap <= 16'b1111111111110000;
		15'h34f4: char_row_bitmap <= 16'b1111111111111000;
		15'h34f5: char_row_bitmap <= 16'b1111111111111100;
		15'h34f6: char_row_bitmap <= 16'b1111111111111110;
		15'h34f7: char_row_bitmap <= 16'b1111111111111111;
		15'h34f8: char_row_bitmap <= 16'b0000000111111111;
		15'h34f9: char_row_bitmap <= 16'b0000001111111111;
		15'h34fa: char_row_bitmap <= 16'b0000011111111111;
		15'h34fb: char_row_bitmap <= 16'b0001111111111111;
		15'h34fc: char_row_bitmap <= 16'b0011111111111111;
		15'h34fd: char_row_bitmap <= 16'b1111111111111111;
		15'h34fe: char_row_bitmap <= 16'b1111111111111111;
		15'h34ff: char_row_bitmap <= 16'b1111111111111111;
		15'h3500: char_row_bitmap <= 16'b1111111111111111;
		15'h3501: char_row_bitmap <= 16'b1111111111111111;
		15'h3502: char_row_bitmap <= 16'b1111111111111111;
		15'h3503: char_row_bitmap <= 16'b1111111111111111;
		15'h3504: char_row_bitmap <= 16'b1111111111111111;
		15'h3505: char_row_bitmap <= 16'b1111111111111111;
		15'h3506: char_row_bitmap <= 16'b1111111111111111;
		15'h3507: char_row_bitmap <= 16'b1111111111111111;
		15'h3508: char_row_bitmap <= 16'b1111111111111111;
		15'h3509: char_row_bitmap <= 16'b1111111111111111;
		15'h350a: char_row_bitmap <= 16'b1111111111111111;
		15'h350b: char_row_bitmap <= 16'b1111111111111111;
		15'h350c: char_row_bitmap <= 16'b0000000000000011;
		15'h350d: char_row_bitmap <= 16'b0000000000001111;
		15'h350e: char_row_bitmap <= 16'b0000000001111111;
		15'h350f: char_row_bitmap <= 16'b0000001111111111;
		15'h3510: char_row_bitmap <= 16'b0000111111111111;
		15'h3511: char_row_bitmap <= 16'b0011111111111111;
		15'h3512: char_row_bitmap <= 16'b1111111111111111;
		15'h3513: char_row_bitmap <= 16'b1111111111111111;
		15'h3514: char_row_bitmap <= 16'b1111111111111111;
		15'h3515: char_row_bitmap <= 16'b1111111111111111;
		15'h3516: char_row_bitmap <= 16'b1111111111111111;
		15'h3517: char_row_bitmap <= 16'b1111111111111111;
		15'h3518: char_row_bitmap <= 16'b1111111111111111;
		15'h3519: char_row_bitmap <= 16'b1111111111111111;
		15'h351a: char_row_bitmap <= 16'b1111111111111111;
		15'h351b: char_row_bitmap <= 16'b1111111111111111;
		15'h351c: char_row_bitmap <= 16'b1111111111111111;
		15'h351d: char_row_bitmap <= 16'b1111111111111111;
		15'h351e: char_row_bitmap <= 16'b1111111111111111;
		15'h351f: char_row_bitmap <= 16'b1111111111111111;
		15'h3520: char_row_bitmap <= 16'b0000000011111111;
		15'h3521: char_row_bitmap <= 16'b0000000111111111;
		15'h3522: char_row_bitmap <= 16'b0000000111111111;
		15'h3523: char_row_bitmap <= 16'b0000001111111111;
		15'h3524: char_row_bitmap <= 16'b0000011111111111;
		15'h3525: char_row_bitmap <= 16'b0000011111111111;
		15'h3526: char_row_bitmap <= 16'b0000111111111111;
		15'h3527: char_row_bitmap <= 16'b0000111111111111;
		15'h3528: char_row_bitmap <= 16'b0001111111111111;
		15'h3529: char_row_bitmap <= 16'b0001111111111111;
		15'h352a: char_row_bitmap <= 16'b0011111111111111;
		15'h352b: char_row_bitmap <= 16'b0111111111111111;
		15'h352c: char_row_bitmap <= 16'b0111111111111111;
		15'h352d: char_row_bitmap <= 16'b1111111111111111;
		15'h352e: char_row_bitmap <= 16'b1111111111111111;
		15'h352f: char_row_bitmap <= 16'b1111111111111111;
		15'h3530: char_row_bitmap <= 16'b1111111111111111;
		15'h3531: char_row_bitmap <= 16'b1111111111111111;
		15'h3532: char_row_bitmap <= 16'b1111111111111111;
		15'h3533: char_row_bitmap <= 16'b1111111111111111;
		15'h3534: char_row_bitmap <= 16'b0000000000000001;
		15'h3535: char_row_bitmap <= 16'b0000000000000011;
		15'h3536: char_row_bitmap <= 16'b0000000000000111;
		15'h3537: char_row_bitmap <= 16'b0000000000001111;
		15'h3538: char_row_bitmap <= 16'b0000000000011111;
		15'h3539: char_row_bitmap <= 16'b0000000000111111;
		15'h353a: char_row_bitmap <= 16'b0000000011111111;
		15'h353b: char_row_bitmap <= 16'b0000000111111111;
		15'h353c: char_row_bitmap <= 16'b0000001111111111;
		15'h353d: char_row_bitmap <= 16'b0000011111111111;
		15'h353e: char_row_bitmap <= 16'b0000111111111111;
		15'h353f: char_row_bitmap <= 16'b0001111111111111;
		15'h3540: char_row_bitmap <= 16'b0011111111111111;
		15'h3541: char_row_bitmap <= 16'b0111111111111111;
		15'h3542: char_row_bitmap <= 16'b1111111111111111;
		15'h3543: char_row_bitmap <= 16'b1111111111111111;
		15'h3544: char_row_bitmap <= 16'b1111111111111111;
		15'h3545: char_row_bitmap <= 16'b1111111111111111;
		15'h3546: char_row_bitmap <= 16'b1111111111111111;
		15'h3547: char_row_bitmap <= 16'b1111111111111111;
		15'h3548: char_row_bitmap <= 16'b0000000011111111;
		15'h3549: char_row_bitmap <= 16'b0000000111111111;
		15'h354a: char_row_bitmap <= 16'b0000000111111111;
		15'h354b: char_row_bitmap <= 16'b0000000111111111;
		15'h354c: char_row_bitmap <= 16'b0000001111111111;
		15'h354d: char_row_bitmap <= 16'b0000001111111111;
		15'h354e: char_row_bitmap <= 16'b0000011111111111;
		15'h354f: char_row_bitmap <= 16'b0000011111111111;
		15'h3550: char_row_bitmap <= 16'b0000011111111111;
		15'h3551: char_row_bitmap <= 16'b0000111111111111;
		15'h3552: char_row_bitmap <= 16'b0000111111111111;
		15'h3553: char_row_bitmap <= 16'b0001111111111111;
		15'h3554: char_row_bitmap <= 16'b0001111111111111;
		15'h3555: char_row_bitmap <= 16'b0001111111111111;
		15'h3556: char_row_bitmap <= 16'b0011111111111111;
		15'h3557: char_row_bitmap <= 16'b0011111111111111;
		15'h3558: char_row_bitmap <= 16'b0111111111111111;
		15'h3559: char_row_bitmap <= 16'b0111111111111111;
		15'h355a: char_row_bitmap <= 16'b0111111111111111;
		15'h355b: char_row_bitmap <= 16'b1111111111111111;
		15'h355c: char_row_bitmap <= 16'b0000000000000000;
		15'h355d: char_row_bitmap <= 16'b0000000000000000;
		15'h355e: char_row_bitmap <= 16'b0000000000000000;
		15'h355f: char_row_bitmap <= 16'b0000000000000000;
		15'h3560: char_row_bitmap <= 16'b0000000000000000;
		15'h3561: char_row_bitmap <= 16'b0000000000000000;
		15'h3562: char_row_bitmap <= 16'b0000000000000001;
		15'h3563: char_row_bitmap <= 16'b0000000000000111;
		15'h3564: char_row_bitmap <= 16'b0000000000011111;
		15'h3565: char_row_bitmap <= 16'b0000000001111111;
		15'h3566: char_row_bitmap <= 16'b0000000111111111;
		15'h3567: char_row_bitmap <= 16'b0000011111111111;
		15'h3568: char_row_bitmap <= 16'b0001111111111111;
		15'h3569: char_row_bitmap <= 16'b0111111111111111;
		15'h356a: char_row_bitmap <= 16'b1111111111111111;
		15'h356b: char_row_bitmap <= 16'b1111111111111111;
		15'h356c: char_row_bitmap <= 16'b1111111111111111;
		15'h356d: char_row_bitmap <= 16'b1111111111111111;
		15'h356e: char_row_bitmap <= 16'b1111111111111111;
		15'h356f: char_row_bitmap <= 16'b1111111111111111;
		15'h3570: char_row_bitmap <= 16'b1111111111111111;
		15'h3571: char_row_bitmap <= 16'b0111111111111111;
		15'h3572: char_row_bitmap <= 16'b0011111111111111;
		15'h3573: char_row_bitmap <= 16'b0001111111111111;
		15'h3574: char_row_bitmap <= 16'b0000111111111111;
		15'h3575: char_row_bitmap <= 16'b0000011111111111;
		15'h3576: char_row_bitmap <= 16'b0000001111111111;
		15'h3577: char_row_bitmap <= 16'b0000000111111111;
		15'h3578: char_row_bitmap <= 16'b0000000011111111;
		15'h3579: char_row_bitmap <= 16'b0000000001111111;
		15'h357a: char_row_bitmap <= 16'b0000000001111111;
		15'h357b: char_row_bitmap <= 16'b0000000011111111;
		15'h357c: char_row_bitmap <= 16'b0000000111111111;
		15'h357d: char_row_bitmap <= 16'b0000001111111111;
		15'h357e: char_row_bitmap <= 16'b0000011111111111;
		15'h357f: char_row_bitmap <= 16'b0000111111111111;
		15'h3580: char_row_bitmap <= 16'b0001111111111111;
		15'h3581: char_row_bitmap <= 16'b0011111111111111;
		15'h3582: char_row_bitmap <= 16'b0111111111111111;
		15'h3583: char_row_bitmap <= 16'b1111111111111111;
		15'h3584: char_row_bitmap <= 16'b1000000000000001;
		15'h3585: char_row_bitmap <= 16'b1100000000000011;
		15'h3586: char_row_bitmap <= 16'b1110000000000111;
		15'h3587: char_row_bitmap <= 16'b1111000000001111;
		15'h3588: char_row_bitmap <= 16'b1111100000011111;
		15'h3589: char_row_bitmap <= 16'b1111110000111111;
		15'h358a: char_row_bitmap <= 16'b1111111001111111;
		15'h358b: char_row_bitmap <= 16'b1111111111111111;
		15'h358c: char_row_bitmap <= 16'b1111111111111111;
		15'h358d: char_row_bitmap <= 16'b1111111111111111;
		15'h358e: char_row_bitmap <= 16'b1111111111111111;
		15'h358f: char_row_bitmap <= 16'b1111111111111111;
		15'h3590: char_row_bitmap <= 16'b1111111111111111;
		15'h3591: char_row_bitmap <= 16'b1111111111111111;
		15'h3592: char_row_bitmap <= 16'b1111111111111111;
		15'h3593: char_row_bitmap <= 16'b1111111111111111;
		15'h3594: char_row_bitmap <= 16'b1111111111111111;
		15'h3595: char_row_bitmap <= 16'b1111111111111111;
		15'h3596: char_row_bitmap <= 16'b1111111111111111;
		15'h3597: char_row_bitmap <= 16'b1111111111111111;
		15'h3598: char_row_bitmap <= 16'b0000000000000000;
		15'h3599: char_row_bitmap <= 16'b0000000000000000;
		15'h359a: char_row_bitmap <= 16'b0000000000000000;
		15'h359b: char_row_bitmap <= 16'b0000000000000000;
		15'h359c: char_row_bitmap <= 16'b0000000000000000;
		15'h359d: char_row_bitmap <= 16'b0000000110000000;
		15'h359e: char_row_bitmap <= 16'b0000000110000000;
		15'h359f: char_row_bitmap <= 16'b0000001111000000;
		15'h35a0: char_row_bitmap <= 16'b0000001111000000;
		15'h35a1: char_row_bitmap <= 16'b0000011111100000;
		15'h35a2: char_row_bitmap <= 16'b0000011111100000;
		15'h35a3: char_row_bitmap <= 16'b0000111111110000;
		15'h35a4: char_row_bitmap <= 16'b0000111111110000;
		15'h35a5: char_row_bitmap <= 16'b0001111111111000;
		15'h35a6: char_row_bitmap <= 16'b0001111111111000;
		15'h35a7: char_row_bitmap <= 16'b0000000000000000;
		15'h35a8: char_row_bitmap <= 16'b0000000000000000;
		15'h35a9: char_row_bitmap <= 16'b0000000000000000;
		15'h35aa: char_row_bitmap <= 16'b0000000000000000;
		15'h35ab: char_row_bitmap <= 16'b0000000000000000;
		15'h35ac: char_row_bitmap <= 16'b0000000000000000;
		15'h35ad: char_row_bitmap <= 16'b0000000000000000;
		15'h35ae: char_row_bitmap <= 16'b0000000000000000;
		15'h35af: char_row_bitmap <= 16'b0000010000000000;
		15'h35b0: char_row_bitmap <= 16'b0000011000000000;
		15'h35b1: char_row_bitmap <= 16'b0000011100000000;
		15'h35b2: char_row_bitmap <= 16'b0000011110000000;
		15'h35b3: char_row_bitmap <= 16'b0000011111000000;
		15'h35b4: char_row_bitmap <= 16'b0000011111100000;
		15'h35b5: char_row_bitmap <= 16'b0000011111110000;
		15'h35b6: char_row_bitmap <= 16'b0000011111110000;
		15'h35b7: char_row_bitmap <= 16'b0000011111100000;
		15'h35b8: char_row_bitmap <= 16'b0000011111000000;
		15'h35b9: char_row_bitmap <= 16'b0000011110000000;
		15'h35ba: char_row_bitmap <= 16'b0000011100000000;
		15'h35bb: char_row_bitmap <= 16'b0000011000000000;
		15'h35bc: char_row_bitmap <= 16'b0000010000000000;
		15'h35bd: char_row_bitmap <= 16'b0000000000000000;
		15'h35be: char_row_bitmap <= 16'b0000000000000000;
		15'h35bf: char_row_bitmap <= 16'b0000000000000000;
		15'h35c0: char_row_bitmap <= 16'b0000000000000000;
		15'h35c1: char_row_bitmap <= 16'b0000000000000000;
		15'h35c2: char_row_bitmap <= 16'b0000000000000000;
		15'h35c3: char_row_bitmap <= 16'b0000000000000000;
		15'h35c4: char_row_bitmap <= 16'b0000000000000000;
		15'h35c5: char_row_bitmap <= 16'b0000000000000000;
		15'h35c6: char_row_bitmap <= 16'b0000000000000000;
		15'h35c7: char_row_bitmap <= 16'b0000000000000000;
		15'h35c8: char_row_bitmap <= 16'b0000000000000000;
		15'h35c9: char_row_bitmap <= 16'b0000000000000000;
		15'h35ca: char_row_bitmap <= 16'b0000000000000000;
		15'h35cb: char_row_bitmap <= 16'b0000000000000000;
		15'h35cc: char_row_bitmap <= 16'b0000000000000000;
		15'h35cd: char_row_bitmap <= 16'b0000000000000000;
		15'h35ce: char_row_bitmap <= 16'b0000000000000001;
		15'h35cf: char_row_bitmap <= 16'b0000000000000011;
		15'h35d0: char_row_bitmap <= 16'b0000000000000111;
		15'h35d1: char_row_bitmap <= 16'b0000000000011111;
		15'h35d2: char_row_bitmap <= 16'b0000000000111111;
		15'h35d3: char_row_bitmap <= 16'b0000000011111111;
		15'h35d4: char_row_bitmap <= 16'b0000000000000000;
		15'h35d5: char_row_bitmap <= 16'b0000000000000000;
		15'h35d6: char_row_bitmap <= 16'b0000000000000000;
		15'h35d7: char_row_bitmap <= 16'b0000000000000000;
		15'h35d8: char_row_bitmap <= 16'b0000000000000000;
		15'h35d9: char_row_bitmap <= 16'b0000000000000000;
		15'h35da: char_row_bitmap <= 16'b0000000000000000;
		15'h35db: char_row_bitmap <= 16'b0000000000000000;
		15'h35dc: char_row_bitmap <= 16'b0000000000000000;
		15'h35dd: char_row_bitmap <= 16'b0000000000000000;
		15'h35de: char_row_bitmap <= 16'b0000000000000000;
		15'h35df: char_row_bitmap <= 16'b0000000000000000;
		15'h35e0: char_row_bitmap <= 16'b0000000000000000;
		15'h35e1: char_row_bitmap <= 16'b0000000000000000;
		15'h35e2: char_row_bitmap <= 16'b0000000000000011;
		15'h35e3: char_row_bitmap <= 16'b0000000000001111;
		15'h35e4: char_row_bitmap <= 16'b0000000001111111;
		15'h35e5: char_row_bitmap <= 16'b0000001111111111;
		15'h35e6: char_row_bitmap <= 16'b0001111111111111;
		15'h35e7: char_row_bitmap <= 16'b0111111111111111;
		15'h35e8: char_row_bitmap <= 16'b0000000000000000;
		15'h35e9: char_row_bitmap <= 16'b0000000000000000;
		15'h35ea: char_row_bitmap <= 16'b0000000000000000;
		15'h35eb: char_row_bitmap <= 16'b0000000000000000;
		15'h35ec: char_row_bitmap <= 16'b0000000000000000;
		15'h35ed: char_row_bitmap <= 16'b0000000000000000;
		15'h35ee: char_row_bitmap <= 16'b0000000000000001;
		15'h35ef: char_row_bitmap <= 16'b0000000000000001;
		15'h35f0: char_row_bitmap <= 16'b0000000000000011;
		15'h35f1: char_row_bitmap <= 16'b0000000000000011;
		15'h35f2: char_row_bitmap <= 16'b0000000000000111;
		15'h35f3: char_row_bitmap <= 16'b0000000000000111;
		15'h35f4: char_row_bitmap <= 16'b0000000000001111;
		15'h35f5: char_row_bitmap <= 16'b0000000000001111;
		15'h35f6: char_row_bitmap <= 16'b0000000000011111;
		15'h35f7: char_row_bitmap <= 16'b0000000000011111;
		15'h35f8: char_row_bitmap <= 16'b0000000000111111;
		15'h35f9: char_row_bitmap <= 16'b0000000001111111;
		15'h35fa: char_row_bitmap <= 16'b0000000001111111;
		15'h35fb: char_row_bitmap <= 16'b0000000011111111;
		15'h35fc: char_row_bitmap <= 16'b0000000000000000;
		15'h35fd: char_row_bitmap <= 16'b0000000000000000;
		15'h35fe: char_row_bitmap <= 16'b0000000000000000;
		15'h35ff: char_row_bitmap <= 16'b0000000000000000;
		15'h3600: char_row_bitmap <= 16'b0000000000000000;
		15'h3601: char_row_bitmap <= 16'b0000000000000000;
		15'h3602: char_row_bitmap <= 16'b0000000000000000;
		15'h3603: char_row_bitmap <= 16'b0000000000000001;
		15'h3604: char_row_bitmap <= 16'b0000000000000011;
		15'h3605: char_row_bitmap <= 16'b0000000000001111;
		15'h3606: char_row_bitmap <= 16'b0000000000011111;
		15'h3607: char_row_bitmap <= 16'b0000000000111111;
		15'h3608: char_row_bitmap <= 16'b0000000001111111;
		15'h3609: char_row_bitmap <= 16'b0000000111111111;
		15'h360a: char_row_bitmap <= 16'b0000001111111111;
		15'h360b: char_row_bitmap <= 16'b0000011111111111;
		15'h360c: char_row_bitmap <= 16'b0000111111111111;
		15'h360d: char_row_bitmap <= 16'b0001111111111111;
		15'h360e: char_row_bitmap <= 16'b0011111111111111;
		15'h360f: char_row_bitmap <= 16'b1111111111111111;
		15'h3610: char_row_bitmap <= 16'b0000000000000001;
		15'h3611: char_row_bitmap <= 16'b0000000000000001;
		15'h3612: char_row_bitmap <= 16'b0000000000000011;
		15'h3613: char_row_bitmap <= 16'b0000000000000011;
		15'h3614: char_row_bitmap <= 16'b0000000000000011;
		15'h3615: char_row_bitmap <= 16'b0000000000000111;
		15'h3616: char_row_bitmap <= 16'b0000000000000111;
		15'h3617: char_row_bitmap <= 16'b0000000000000111;
		15'h3618: char_row_bitmap <= 16'b0000000000001111;
		15'h3619: char_row_bitmap <= 16'b0000000000001111;
		15'h361a: char_row_bitmap <= 16'b0000000000001111;
		15'h361b: char_row_bitmap <= 16'b0000000000011111;
		15'h361c: char_row_bitmap <= 16'b0000000000011111;
		15'h361d: char_row_bitmap <= 16'b0000000000011111;
		15'h361e: char_row_bitmap <= 16'b0000000000111111;
		15'h361f: char_row_bitmap <= 16'b0000000000111111;
		15'h3620: char_row_bitmap <= 16'b0000000001111111;
		15'h3621: char_row_bitmap <= 16'b0000000001111111;
		15'h3622: char_row_bitmap <= 16'b0000000001111111;
		15'h3623: char_row_bitmap <= 16'b0000000011111111;
		15'h3624: char_row_bitmap <= 16'b0000000000000001;
		15'h3625: char_row_bitmap <= 16'b0000000000000011;
		15'h3626: char_row_bitmap <= 16'b0000000000000011;
		15'h3627: char_row_bitmap <= 16'b0000000000000111;
		15'h3628: char_row_bitmap <= 16'b0000000000001111;
		15'h3629: char_row_bitmap <= 16'b0000000000001111;
		15'h362a: char_row_bitmap <= 16'b0000000000011111;
		15'h362b: char_row_bitmap <= 16'b0000000000111111;
		15'h362c: char_row_bitmap <= 16'b0000000001111111;
		15'h362d: char_row_bitmap <= 16'b0000000011111111;
		15'h362e: char_row_bitmap <= 16'b0000000011111111;
		15'h362f: char_row_bitmap <= 16'b0000000111111111;
		15'h3630: char_row_bitmap <= 16'b0000001111111111;
		15'h3631: char_row_bitmap <= 16'b0000011111111111;
		15'h3632: char_row_bitmap <= 16'b0000111111111111;
		15'h3633: char_row_bitmap <= 16'b0000111111111111;
		15'h3634: char_row_bitmap <= 16'b0001111111111111;
		15'h3635: char_row_bitmap <= 16'b0011111111111111;
		15'h3636: char_row_bitmap <= 16'b0111111111111111;
		15'h3637: char_row_bitmap <= 16'b1111111111111111;
		15'h3638: char_row_bitmap <= 16'b1111111110000000;
		15'h3639: char_row_bitmap <= 16'b1111111111000000;
		15'h363a: char_row_bitmap <= 16'b1111111111100000;
		15'h363b: char_row_bitmap <= 16'b1111111111111000;
		15'h363c: char_row_bitmap <= 16'b1111111111111100;
		15'h363d: char_row_bitmap <= 16'b1111111111111111;
		15'h363e: char_row_bitmap <= 16'b1111111111111111;
		15'h363f: char_row_bitmap <= 16'b1111111111111111;
		15'h3640: char_row_bitmap <= 16'b1111111111111111;
		15'h3641: char_row_bitmap <= 16'b1111111111111111;
		15'h3642: char_row_bitmap <= 16'b1111111111111111;
		15'h3643: char_row_bitmap <= 16'b1111111111111111;
		15'h3644: char_row_bitmap <= 16'b1111111111111111;
		15'h3645: char_row_bitmap <= 16'b1111111111111111;
		15'h3646: char_row_bitmap <= 16'b1111111111111111;
		15'h3647: char_row_bitmap <= 16'b1111111111111111;
		15'h3648: char_row_bitmap <= 16'b1111111111111111;
		15'h3649: char_row_bitmap <= 16'b1111111111111111;
		15'h364a: char_row_bitmap <= 16'b1111111111111111;
		15'h364b: char_row_bitmap <= 16'b1111111111111111;
		15'h364c: char_row_bitmap <= 16'b1100000000000000;
		15'h364d: char_row_bitmap <= 16'b1111000000000000;
		15'h364e: char_row_bitmap <= 16'b1111111000000000;
		15'h364f: char_row_bitmap <= 16'b1111111111000000;
		15'h3650: char_row_bitmap <= 16'b1111111111110000;
		15'h3651: char_row_bitmap <= 16'b1111111111111100;
		15'h3652: char_row_bitmap <= 16'b1111111111111111;
		15'h3653: char_row_bitmap <= 16'b1111111111111111;
		15'h3654: char_row_bitmap <= 16'b1111111111111111;
		15'h3655: char_row_bitmap <= 16'b1111111111111111;
		15'h3656: char_row_bitmap <= 16'b1111111111111111;
		15'h3657: char_row_bitmap <= 16'b1111111111111111;
		15'h3658: char_row_bitmap <= 16'b1111111111111111;
		15'h3659: char_row_bitmap <= 16'b1111111111111111;
		15'h365a: char_row_bitmap <= 16'b1111111111111111;
		15'h365b: char_row_bitmap <= 16'b1111111111111111;
		15'h365c: char_row_bitmap <= 16'b1111111111111111;
		15'h365d: char_row_bitmap <= 16'b1111111111111111;
		15'h365e: char_row_bitmap <= 16'b1111111111111111;
		15'h365f: char_row_bitmap <= 16'b1111111111111111;
		15'h3660: char_row_bitmap <= 16'b1111111100000000;
		15'h3661: char_row_bitmap <= 16'b1111111110000000;
		15'h3662: char_row_bitmap <= 16'b1111111110000000;
		15'h3663: char_row_bitmap <= 16'b1111111111000000;
		15'h3664: char_row_bitmap <= 16'b1111111111100000;
		15'h3665: char_row_bitmap <= 16'b1111111111100000;
		15'h3666: char_row_bitmap <= 16'b1111111111110000;
		15'h3667: char_row_bitmap <= 16'b1111111111110000;
		15'h3668: char_row_bitmap <= 16'b1111111111111000;
		15'h3669: char_row_bitmap <= 16'b1111111111111000;
		15'h366a: char_row_bitmap <= 16'b1111111111111100;
		15'h366b: char_row_bitmap <= 16'b1111111111111110;
		15'h366c: char_row_bitmap <= 16'b1111111111111110;
		15'h366d: char_row_bitmap <= 16'b1111111111111111;
		15'h366e: char_row_bitmap <= 16'b1111111111111111;
		15'h366f: char_row_bitmap <= 16'b1111111111111111;
		15'h3670: char_row_bitmap <= 16'b1111111111111111;
		15'h3671: char_row_bitmap <= 16'b1111111111111111;
		15'h3672: char_row_bitmap <= 16'b1111111111111111;
		15'h3673: char_row_bitmap <= 16'b1111111111111111;
		15'h3674: char_row_bitmap <= 16'b1000000000000000;
		15'h3675: char_row_bitmap <= 16'b1100000000000000;
		15'h3676: char_row_bitmap <= 16'b1110000000000000;
		15'h3677: char_row_bitmap <= 16'b1111000000000000;
		15'h3678: char_row_bitmap <= 16'b1111100000000000;
		15'h3679: char_row_bitmap <= 16'b1111110000000000;
		15'h367a: char_row_bitmap <= 16'b1111111100000000;
		15'h367b: char_row_bitmap <= 16'b1111111110000000;
		15'h367c: char_row_bitmap <= 16'b1111111111000000;
		15'h367d: char_row_bitmap <= 16'b1111111111100000;
		15'h367e: char_row_bitmap <= 16'b1111111111110000;
		15'h367f: char_row_bitmap <= 16'b1111111111111000;
		15'h3680: char_row_bitmap <= 16'b1111111111111100;
		15'h3681: char_row_bitmap <= 16'b1111111111111110;
		15'h3682: char_row_bitmap <= 16'b1111111111111111;
		15'h3683: char_row_bitmap <= 16'b1111111111111111;
		15'h3684: char_row_bitmap <= 16'b1111111111111111;
		15'h3685: char_row_bitmap <= 16'b1111111111111111;
		15'h3686: char_row_bitmap <= 16'b1111111111111111;
		15'h3687: char_row_bitmap <= 16'b1111111111111111;
		15'h3688: char_row_bitmap <= 16'b1111111100000000;
		15'h3689: char_row_bitmap <= 16'b1111111110000000;
		15'h368a: char_row_bitmap <= 16'b1111111110000000;
		15'h368b: char_row_bitmap <= 16'b1111111110000000;
		15'h368c: char_row_bitmap <= 16'b1111111111000000;
		15'h368d: char_row_bitmap <= 16'b1111111111000000;
		15'h368e: char_row_bitmap <= 16'b1111111111100000;
		15'h368f: char_row_bitmap <= 16'b1111111111100000;
		15'h3690: char_row_bitmap <= 16'b1111111111100000;
		15'h3691: char_row_bitmap <= 16'b1111111111110000;
		15'h3692: char_row_bitmap <= 16'b1111111111110000;
		15'h3693: char_row_bitmap <= 16'b1111111111111000;
		15'h3694: char_row_bitmap <= 16'b1111111111111000;
		15'h3695: char_row_bitmap <= 16'b1111111111111000;
		15'h3696: char_row_bitmap <= 16'b1111111111111100;
		15'h3697: char_row_bitmap <= 16'b1111111111111100;
		15'h3698: char_row_bitmap <= 16'b1111111111111110;
		15'h3699: char_row_bitmap <= 16'b1111111111111110;
		15'h369a: char_row_bitmap <= 16'b1111111111111110;
		15'h369b: char_row_bitmap <= 16'b1111111111111111;
		15'h369c: char_row_bitmap <= 16'b0000000000000000;
		15'h369d: char_row_bitmap <= 16'b0000000000000000;
		15'h369e: char_row_bitmap <= 16'b0000000000000000;
		15'h369f: char_row_bitmap <= 16'b0000000000000000;
		15'h36a0: char_row_bitmap <= 16'b0000000000000000;
		15'h36a1: char_row_bitmap <= 16'b0000000000000000;
		15'h36a2: char_row_bitmap <= 16'b1000000000000000;
		15'h36a3: char_row_bitmap <= 16'b1110000000000000;
		15'h36a4: char_row_bitmap <= 16'b1111100000000000;
		15'h36a5: char_row_bitmap <= 16'b1111111000000000;
		15'h36a6: char_row_bitmap <= 16'b1111111110000000;
		15'h36a7: char_row_bitmap <= 16'b1111111111100000;
		15'h36a8: char_row_bitmap <= 16'b1111111111111000;
		15'h36a9: char_row_bitmap <= 16'b1111111111111110;
		15'h36aa: char_row_bitmap <= 16'b1111111111111111;
		15'h36ab: char_row_bitmap <= 16'b1111111111111111;
		15'h36ac: char_row_bitmap <= 16'b1111111111111111;
		15'h36ad: char_row_bitmap <= 16'b1111111111111111;
		15'h36ae: char_row_bitmap <= 16'b1111111111111111;
		15'h36af: char_row_bitmap <= 16'b1111111111111111;
		15'h36b0: char_row_bitmap <= 16'b1111111111111111;
		15'h36b1: char_row_bitmap <= 16'b1111111111111110;
		15'h36b2: char_row_bitmap <= 16'b1111111111111100;
		15'h36b3: char_row_bitmap <= 16'b1111111111111000;
		15'h36b4: char_row_bitmap <= 16'b1111111111110000;
		15'h36b5: char_row_bitmap <= 16'b1111111111100000;
		15'h36b6: char_row_bitmap <= 16'b1111111111000000;
		15'h36b7: char_row_bitmap <= 16'b1111111110000000;
		15'h36b8: char_row_bitmap <= 16'b1111111100000000;
		15'h36b9: char_row_bitmap <= 16'b1111111000000000;
		15'h36ba: char_row_bitmap <= 16'b1111111000000000;
		15'h36bb: char_row_bitmap <= 16'b1111111100000000;
		15'h36bc: char_row_bitmap <= 16'b1111111110000000;
		15'h36bd: char_row_bitmap <= 16'b1111111111000000;
		15'h36be: char_row_bitmap <= 16'b1111111111100000;
		15'h36bf: char_row_bitmap <= 16'b1111111111110000;
		15'h36c0: char_row_bitmap <= 16'b1111111111111000;
		15'h36c1: char_row_bitmap <= 16'b1111111111111100;
		15'h36c2: char_row_bitmap <= 16'b1111111111111110;
		15'h36c3: char_row_bitmap <= 16'b1111111111111111;
		15'h36c4: char_row_bitmap <= 16'b1111111111111111;
		15'h36c5: char_row_bitmap <= 16'b1111111111111111;
		15'h36c6: char_row_bitmap <= 16'b1111111111111111;
		15'h36c7: char_row_bitmap <= 16'b1111111111111111;
		15'h36c8: char_row_bitmap <= 16'b1111111111111111;
		15'h36c9: char_row_bitmap <= 16'b1111111111111111;
		15'h36ca: char_row_bitmap <= 16'b1111111111111111;
		15'h36cb: char_row_bitmap <= 16'b1111111111111111;
		15'h36cc: char_row_bitmap <= 16'b1111111111111111;
		15'h36cd: char_row_bitmap <= 16'b1111111111111111;
		15'h36ce: char_row_bitmap <= 16'b1111111111111111;
		15'h36cf: char_row_bitmap <= 16'b1111111111111111;
		15'h36d0: char_row_bitmap <= 16'b1111111111111111;
		15'h36d1: char_row_bitmap <= 16'b1111111001111111;
		15'h36d2: char_row_bitmap <= 16'b1111110000111111;
		15'h36d3: char_row_bitmap <= 16'b1111100000011111;
		15'h36d4: char_row_bitmap <= 16'b1111000000001111;
		15'h36d5: char_row_bitmap <= 16'b1110000000000111;
		15'h36d6: char_row_bitmap <= 16'b1100000000000011;
		15'h36d7: char_row_bitmap <= 16'b1000000000000001;
		15'h36d8: char_row_bitmap <= 16'b0000000000000000;
		15'h36d9: char_row_bitmap <= 16'b0000000000000000;
		15'h36da: char_row_bitmap <= 16'b0000000000000000;
		15'h36db: char_row_bitmap <= 16'b0000000000000000;
		15'h36dc: char_row_bitmap <= 16'b0000000000000000;
		15'h36dd: char_row_bitmap <= 16'b0001111111111000;
		15'h36de: char_row_bitmap <= 16'b0001111111111000;
		15'h36df: char_row_bitmap <= 16'b0000111111110000;
		15'h36e0: char_row_bitmap <= 16'b0000111111110000;
		15'h36e1: char_row_bitmap <= 16'b0000011111100000;
		15'h36e2: char_row_bitmap <= 16'b0000011111100000;
		15'h36e3: char_row_bitmap <= 16'b0000001111000000;
		15'h36e4: char_row_bitmap <= 16'b0000001111000000;
		15'h36e5: char_row_bitmap <= 16'b0000000110000000;
		15'h36e6: char_row_bitmap <= 16'b0000000110000000;
		15'h36e7: char_row_bitmap <= 16'b0000000000000000;
		15'h36e8: char_row_bitmap <= 16'b0000000000000000;
		15'h36e9: char_row_bitmap <= 16'b0000000000000000;
		15'h36ea: char_row_bitmap <= 16'b0000000000000000;
		15'h36eb: char_row_bitmap <= 16'b0000000000000000;
		15'h36ec: char_row_bitmap <= 16'b0000000000000000;
		15'h36ed: char_row_bitmap <= 16'b0000000000000000;
		15'h36ee: char_row_bitmap <= 16'b0000000000000000;
		15'h36ef: char_row_bitmap <= 16'b0000000000100000;
		15'h36f0: char_row_bitmap <= 16'b0000000001100000;
		15'h36f1: char_row_bitmap <= 16'b0000000011100000;
		15'h36f2: char_row_bitmap <= 16'b0000000111100000;
		15'h36f3: char_row_bitmap <= 16'b0000001111100000;
		15'h36f4: char_row_bitmap <= 16'b0000011111100000;
		15'h36f5: char_row_bitmap <= 16'b0000111111100000;
		15'h36f6: char_row_bitmap <= 16'b0000111111100000;
		15'h36f7: char_row_bitmap <= 16'b0000011111100000;
		15'h36f8: char_row_bitmap <= 16'b0000001111100000;
		15'h36f9: char_row_bitmap <= 16'b0000000111100000;
		15'h36fa: char_row_bitmap <= 16'b0000000011100000;
		15'h36fb: char_row_bitmap <= 16'b0000000001100000;
		15'h36fc: char_row_bitmap <= 16'b0000000000100000;
		15'h36fd: char_row_bitmap <= 16'b0000000000000000;
		15'h36fe: char_row_bitmap <= 16'b0000000000000000;
		15'h36ff: char_row_bitmap <= 16'b0000000000000000;
		15'h3700: char_row_bitmap <= 16'b1111111111111111;
		15'h3701: char_row_bitmap <= 16'b1111111111111111;
		15'h3702: char_row_bitmap <= 16'b1111111111111111;
		15'h3703: char_row_bitmap <= 16'b1111111111111111;
		15'h3704: char_row_bitmap <= 16'b1111111111111111;
		15'h3705: char_row_bitmap <= 16'b1111111111111111;
		15'h3706: char_row_bitmap <= 16'b1111111111111111;
		15'h3707: char_row_bitmap <= 16'b1111111111111111;
		15'h3708: char_row_bitmap <= 16'b1111111111111111;
		15'h3709: char_row_bitmap <= 16'b1111111111111111;
		15'h370a: char_row_bitmap <= 16'b1111111111111111;
		15'h370b: char_row_bitmap <= 16'b1111111111111111;
		15'h370c: char_row_bitmap <= 16'b1111111111111111;
		15'h370d: char_row_bitmap <= 16'b1111111111111111;
		15'h370e: char_row_bitmap <= 16'b1111111111111111;
		15'h370f: char_row_bitmap <= 16'b0011111111111111;
		15'h3710: char_row_bitmap <= 16'b0001111111111111;
		15'h3711: char_row_bitmap <= 16'b0000011111111111;
		15'h3712: char_row_bitmap <= 16'b0000001111111111;
		15'h3713: char_row_bitmap <= 16'b0000000111111111;
		15'h3714: char_row_bitmap <= 16'b1111111111111111;
		15'h3715: char_row_bitmap <= 16'b1111111111111111;
		15'h3716: char_row_bitmap <= 16'b1111111111111111;
		15'h3717: char_row_bitmap <= 16'b1111111111111111;
		15'h3718: char_row_bitmap <= 16'b1111111111111111;
		15'h3719: char_row_bitmap <= 16'b1111111111111111;
		15'h371a: char_row_bitmap <= 16'b1111111111111111;
		15'h371b: char_row_bitmap <= 16'b1111111111111111;
		15'h371c: char_row_bitmap <= 16'b1111111111111111;
		15'h371d: char_row_bitmap <= 16'b1111111111111111;
		15'h371e: char_row_bitmap <= 16'b1111111111111111;
		15'h371f: char_row_bitmap <= 16'b1111111111111111;
		15'h3720: char_row_bitmap <= 16'b1111111111111111;
		15'h3721: char_row_bitmap <= 16'b1111111111111111;
		15'h3722: char_row_bitmap <= 16'b0011111111111111;
		15'h3723: char_row_bitmap <= 16'b0000111111111111;
		15'h3724: char_row_bitmap <= 16'b0000001111111111;
		15'h3725: char_row_bitmap <= 16'b0000000001111111;
		15'h3726: char_row_bitmap <= 16'b0000000000001111;
		15'h3727: char_row_bitmap <= 16'b0000000000000011;
		15'h3728: char_row_bitmap <= 16'b1111111111111111;
		15'h3729: char_row_bitmap <= 16'b1111111111111111;
		15'h372a: char_row_bitmap <= 16'b1111111111111111;
		15'h372b: char_row_bitmap <= 16'b1111111111111111;
		15'h372c: char_row_bitmap <= 16'b1111111111111111;
		15'h372d: char_row_bitmap <= 16'b1111111111111111;
		15'h372e: char_row_bitmap <= 16'b1111111111111111;
		15'h372f: char_row_bitmap <= 16'b0111111111111111;
		15'h3730: char_row_bitmap <= 16'b0111111111111111;
		15'h3731: char_row_bitmap <= 16'b0011111111111111;
		15'h3732: char_row_bitmap <= 16'b0001111111111111;
		15'h3733: char_row_bitmap <= 16'b0001111111111111;
		15'h3734: char_row_bitmap <= 16'b0000111111111111;
		15'h3735: char_row_bitmap <= 16'b0000111111111111;
		15'h3736: char_row_bitmap <= 16'b0000011111111111;
		15'h3737: char_row_bitmap <= 16'b0000011111111111;
		15'h3738: char_row_bitmap <= 16'b0000001111111111;
		15'h3739: char_row_bitmap <= 16'b0000000111111111;
		15'h373a: char_row_bitmap <= 16'b0000000111111111;
		15'h373b: char_row_bitmap <= 16'b0000000011111111;
		15'h373c: char_row_bitmap <= 16'b1111111111111111;
		15'h373d: char_row_bitmap <= 16'b0011111111111111;
		15'h373e: char_row_bitmap <= 16'b0001111111111111;
		15'h373f: char_row_bitmap <= 16'b0000111111111111;
		15'h3740: char_row_bitmap <= 16'b0000011111111111;
		15'h3741: char_row_bitmap <= 16'b0000001111111111;
		15'h3742: char_row_bitmap <= 16'b0000000111111111;
		15'h3743: char_row_bitmap <= 16'b0000000001111111;
		15'h3744: char_row_bitmap <= 16'b0000000000111111;
		15'h3745: char_row_bitmap <= 16'b0000000000011111;
		15'h3746: char_row_bitmap <= 16'b0000000000001111;
		15'h3747: char_row_bitmap <= 16'b0000000000000011;
		15'h3748: char_row_bitmap <= 16'b0000000000000001;
		15'h3749: char_row_bitmap <= 16'b0000000000000000;
		15'h374a: char_row_bitmap <= 16'b0000000000000000;
		15'h374b: char_row_bitmap <= 16'b0000000000000000;
		15'h374c: char_row_bitmap <= 16'b0000000000000000;
		15'h374d: char_row_bitmap <= 16'b0000000000000000;
		15'h374e: char_row_bitmap <= 16'b0000000000000000;
		15'h374f: char_row_bitmap <= 16'b0000000000000000;
		15'h3750: char_row_bitmap <= 16'b1111111111111111;
		15'h3751: char_row_bitmap <= 16'b0111111111111111;
		15'h3752: char_row_bitmap <= 16'b0111111111111111;
		15'h3753: char_row_bitmap <= 16'b0111111111111111;
		15'h3754: char_row_bitmap <= 16'b0011111111111111;
		15'h3755: char_row_bitmap <= 16'b0011111111111111;
		15'h3756: char_row_bitmap <= 16'b0001111111111111;
		15'h3757: char_row_bitmap <= 16'b0001111111111111;
		15'h3758: char_row_bitmap <= 16'b0001111111111111;
		15'h3759: char_row_bitmap <= 16'b0000111111111111;
		15'h375a: char_row_bitmap <= 16'b0000111111111111;
		15'h375b: char_row_bitmap <= 16'b0000011111111111;
		15'h375c: char_row_bitmap <= 16'b0000011111111111;
		15'h375d: char_row_bitmap <= 16'b0000011111111111;
		15'h375e: char_row_bitmap <= 16'b0000001111111111;
		15'h375f: char_row_bitmap <= 16'b0000001111111111;
		15'h3760: char_row_bitmap <= 16'b0000000111111111;
		15'h3761: char_row_bitmap <= 16'b0000000111111111;
		15'h3762: char_row_bitmap <= 16'b0000000111111111;
		15'h3763: char_row_bitmap <= 16'b0000000011111111;
		15'h3764: char_row_bitmap <= 16'b1111111111111111;
		15'h3765: char_row_bitmap <= 16'b0111111111111111;
		15'h3766: char_row_bitmap <= 16'b0011111111111111;
		15'h3767: char_row_bitmap <= 16'b0001111111111111;
		15'h3768: char_row_bitmap <= 16'b0000111111111111;
		15'h3769: char_row_bitmap <= 16'b0000111111111111;
		15'h376a: char_row_bitmap <= 16'b0000011111111111;
		15'h376b: char_row_bitmap <= 16'b0000001111111111;
		15'h376c: char_row_bitmap <= 16'b0000000111111111;
		15'h376d: char_row_bitmap <= 16'b0000000011111111;
		15'h376e: char_row_bitmap <= 16'b0000000011111111;
		15'h376f: char_row_bitmap <= 16'b0000000001111111;
		15'h3770: char_row_bitmap <= 16'b0000000000111111;
		15'h3771: char_row_bitmap <= 16'b0000000000011111;
		15'h3772: char_row_bitmap <= 16'b0000000000001111;
		15'h3773: char_row_bitmap <= 16'b0000000000001111;
		15'h3774: char_row_bitmap <= 16'b0000000000000111;
		15'h3775: char_row_bitmap <= 16'b0000000000000011;
		15'h3776: char_row_bitmap <= 16'b0000000000000011;
		15'h3777: char_row_bitmap <= 16'b0000000000000001;
		15'h3778: char_row_bitmap <= 16'b1111111100000000;
		15'h3779: char_row_bitmap <= 16'b1111110000000000;
		15'h377a: char_row_bitmap <= 16'b1111100000000000;
		15'h377b: char_row_bitmap <= 16'b1110000000000000;
		15'h377c: char_row_bitmap <= 16'b1100000000000000;
		15'h377d: char_row_bitmap <= 16'b1000000000000000;
		15'h377e: char_row_bitmap <= 16'b0000000000000000;
		15'h377f: char_row_bitmap <= 16'b0000000000000000;
		15'h3780: char_row_bitmap <= 16'b0000000000000000;
		15'h3781: char_row_bitmap <= 16'b0000000000000000;
		15'h3782: char_row_bitmap <= 16'b0000000000000000;
		15'h3783: char_row_bitmap <= 16'b0000000000000000;
		15'h3784: char_row_bitmap <= 16'b0000000000000000;
		15'h3785: char_row_bitmap <= 16'b0000000000000000;
		15'h3786: char_row_bitmap <= 16'b0000000000000000;
		15'h3787: char_row_bitmap <= 16'b0000000000000000;
		15'h3788: char_row_bitmap <= 16'b0000000000000000;
		15'h3789: char_row_bitmap <= 16'b0000000000000000;
		15'h378a: char_row_bitmap <= 16'b0000000000000000;
		15'h378b: char_row_bitmap <= 16'b0000000000000000;
		15'h378c: char_row_bitmap <= 16'b1111111111111110;
		15'h378d: char_row_bitmap <= 16'b1111111111111000;
		15'h378e: char_row_bitmap <= 16'b1111111111000000;
		15'h378f: char_row_bitmap <= 16'b1111111000000000;
		15'h3790: char_row_bitmap <= 16'b1111000000000000;
		15'h3791: char_row_bitmap <= 16'b1100000000000000;
		15'h3792: char_row_bitmap <= 16'b0000000000000000;
		15'h3793: char_row_bitmap <= 16'b0000000000000000;
		15'h3794: char_row_bitmap <= 16'b0000000000000000;
		15'h3795: char_row_bitmap <= 16'b0000000000000000;
		15'h3796: char_row_bitmap <= 16'b0000000000000000;
		15'h3797: char_row_bitmap <= 16'b0000000000000000;
		15'h3798: char_row_bitmap <= 16'b0000000000000000;
		15'h3799: char_row_bitmap <= 16'b0000000000000000;
		15'h379a: char_row_bitmap <= 16'b0000000000000000;
		15'h379b: char_row_bitmap <= 16'b0000000000000000;
		15'h379c: char_row_bitmap <= 16'b0000000000000000;
		15'h379d: char_row_bitmap <= 16'b0000000000000000;
		15'h379e: char_row_bitmap <= 16'b0000000000000000;
		15'h379f: char_row_bitmap <= 16'b0000000000000000;
		15'h37a0: char_row_bitmap <= 16'b1111111100000000;
		15'h37a1: char_row_bitmap <= 16'b1111111000000000;
		15'h37a2: char_row_bitmap <= 16'b1111111000000000;
		15'h37a3: char_row_bitmap <= 16'b1111110000000000;
		15'h37a4: char_row_bitmap <= 16'b1111100000000000;
		15'h37a5: char_row_bitmap <= 16'b1111100000000000;
		15'h37a6: char_row_bitmap <= 16'b1111000000000000;
		15'h37a7: char_row_bitmap <= 16'b1111000000000000;
		15'h37a8: char_row_bitmap <= 16'b1110000000000000;
		15'h37a9: char_row_bitmap <= 16'b1110000000000000;
		15'h37aa: char_row_bitmap <= 16'b1100000000000000;
		15'h37ab: char_row_bitmap <= 16'b1100000000000000;
		15'h37ac: char_row_bitmap <= 16'b1000000000000000;
		15'h37ad: char_row_bitmap <= 16'b1000000000000000;
		15'h37ae: char_row_bitmap <= 16'b0000000000000000;
		15'h37af: char_row_bitmap <= 16'b0000000000000000;
		15'h37b0: char_row_bitmap <= 16'b0000000000000000;
		15'h37b1: char_row_bitmap <= 16'b0000000000000000;
		15'h37b2: char_row_bitmap <= 16'b0000000000000000;
		15'h37b3: char_row_bitmap <= 16'b0000000000000000;
		15'h37b4: char_row_bitmap <= 16'b1111111111111110;
		15'h37b5: char_row_bitmap <= 16'b1111111111111100;
		15'h37b6: char_row_bitmap <= 16'b1111111111111000;
		15'h37b7: char_row_bitmap <= 16'b1111111111110000;
		15'h37b8: char_row_bitmap <= 16'b1111111111100000;
		15'h37b9: char_row_bitmap <= 16'b1111111111000000;
		15'h37ba: char_row_bitmap <= 16'b1111111110000000;
		15'h37bb: char_row_bitmap <= 16'b1111111000000000;
		15'h37bc: char_row_bitmap <= 16'b1111110000000000;
		15'h37bd: char_row_bitmap <= 16'b1111100000000000;
		15'h37be: char_row_bitmap <= 16'b1111000000000000;
		15'h37bf: char_row_bitmap <= 16'b1100000000000000;
		15'h37c0: char_row_bitmap <= 16'b1000000000000000;
		15'h37c1: char_row_bitmap <= 16'b0000000000000000;
		15'h37c2: char_row_bitmap <= 16'b0000000000000000;
		15'h37c3: char_row_bitmap <= 16'b0000000000000000;
		15'h37c4: char_row_bitmap <= 16'b0000000000000000;
		15'h37c5: char_row_bitmap <= 16'b0000000000000000;
		15'h37c6: char_row_bitmap <= 16'b0000000000000000;
		15'h37c7: char_row_bitmap <= 16'b0000000000000000;
		15'h37c8: char_row_bitmap <= 16'b1111111100000000;
		15'h37c9: char_row_bitmap <= 16'b1111111000000000;
		15'h37ca: char_row_bitmap <= 16'b1111111000000000;
		15'h37cb: char_row_bitmap <= 16'b1111111000000000;
		15'h37cc: char_row_bitmap <= 16'b1111110000000000;
		15'h37cd: char_row_bitmap <= 16'b1111110000000000;
		15'h37ce: char_row_bitmap <= 16'b1111100000000000;
		15'h37cf: char_row_bitmap <= 16'b1111100000000000;
		15'h37d0: char_row_bitmap <= 16'b1111100000000000;
		15'h37d1: char_row_bitmap <= 16'b1111000000000000;
		15'h37d2: char_row_bitmap <= 16'b1111000000000000;
		15'h37d3: char_row_bitmap <= 16'b1111000000000000;
		15'h37d4: char_row_bitmap <= 16'b1110000000000000;
		15'h37d5: char_row_bitmap <= 16'b1110000000000000;
		15'h37d6: char_row_bitmap <= 16'b1110000000000000;
		15'h37d7: char_row_bitmap <= 16'b1100000000000000;
		15'h37d8: char_row_bitmap <= 16'b1100000000000000;
		15'h37d9: char_row_bitmap <= 16'b1100000000000000;
		15'h37da: char_row_bitmap <= 16'b1000000000000000;
		15'h37db: char_row_bitmap <= 16'b1000000000000000;
		15'h37dc: char_row_bitmap <= 16'b1111111111111111;
		15'h37dd: char_row_bitmap <= 16'b1111111111111111;
		15'h37de: char_row_bitmap <= 16'b1111111111111111;
		15'h37df: char_row_bitmap <= 16'b1111111111111111;
		15'h37e0: char_row_bitmap <= 16'b1111111111111111;
		15'h37e1: char_row_bitmap <= 16'b1111111111111111;
		15'h37e2: char_row_bitmap <= 16'b1111111111111110;
		15'h37e3: char_row_bitmap <= 16'b1111111111111000;
		15'h37e4: char_row_bitmap <= 16'b1111111111100000;
		15'h37e5: char_row_bitmap <= 16'b1111111110000000;
		15'h37e6: char_row_bitmap <= 16'b1111111000000000;
		15'h37e7: char_row_bitmap <= 16'b1111100000000000;
		15'h37e8: char_row_bitmap <= 16'b1110000000000000;
		15'h37e9: char_row_bitmap <= 16'b1000000000000000;
		15'h37ea: char_row_bitmap <= 16'b0000000000000000;
		15'h37eb: char_row_bitmap <= 16'b0000000000000000;
		15'h37ec: char_row_bitmap <= 16'b0000000000000000;
		15'h37ed: char_row_bitmap <= 16'b0000000000000000;
		15'h37ee: char_row_bitmap <= 16'b0000000000000000;
		15'h37ef: char_row_bitmap <= 16'b0000000000000000;
		15'h37f0: char_row_bitmap <= 16'b0000000000000000;
		15'h37f1: char_row_bitmap <= 16'b1000000000000000;
		15'h37f2: char_row_bitmap <= 16'b1100000000000000;
		15'h37f3: char_row_bitmap <= 16'b1110000000000000;
		15'h37f4: char_row_bitmap <= 16'b1111000000000000;
		15'h37f5: char_row_bitmap <= 16'b1111100000000000;
		15'h37f6: char_row_bitmap <= 16'b1111110000000000;
		15'h37f7: char_row_bitmap <= 16'b1111111000000000;
		15'h37f8: char_row_bitmap <= 16'b1111111100000000;
		15'h37f9: char_row_bitmap <= 16'b1111111110000000;
		15'h37fa: char_row_bitmap <= 16'b1111111110000000;
		15'h37fb: char_row_bitmap <= 16'b1111111100000000;
		15'h37fc: char_row_bitmap <= 16'b1111111000000000;
		15'h37fd: char_row_bitmap <= 16'b1111110000000000;
		15'h37fe: char_row_bitmap <= 16'b1111100000000000;
		15'h37ff: char_row_bitmap <= 16'b1111000000000000;
		15'h3800: char_row_bitmap <= 16'b1110000000000000;
		15'h3801: char_row_bitmap <= 16'b1100000000000000;
		15'h3802: char_row_bitmap <= 16'b1000000000000000;
		15'h3803: char_row_bitmap <= 16'b0000000000000000;
		15'h3804: char_row_bitmap <= 16'b0111111111111110;
		15'h3805: char_row_bitmap <= 16'b0011111111111100;
		15'h3806: char_row_bitmap <= 16'b0001111111111000;
		15'h3807: char_row_bitmap <= 16'b0000111111110000;
		15'h3808: char_row_bitmap <= 16'b0000011111100000;
		15'h3809: char_row_bitmap <= 16'b0000001111000000;
		15'h380a: char_row_bitmap <= 16'b0000000110000000;
		15'h380b: char_row_bitmap <= 16'b0000000000000000;
		15'h380c: char_row_bitmap <= 16'b0000000000000000;
		15'h380d: char_row_bitmap <= 16'b0000000000000000;
		15'h380e: char_row_bitmap <= 16'b0000000000000000;
		15'h380f: char_row_bitmap <= 16'b0000000000000000;
		15'h3810: char_row_bitmap <= 16'b0000000000000000;
		15'h3811: char_row_bitmap <= 16'b0000000000000000;
		15'h3812: char_row_bitmap <= 16'b0000000000000000;
		15'h3813: char_row_bitmap <= 16'b0000000000000000;
		15'h3814: char_row_bitmap <= 16'b0000000000000000;
		15'h3815: char_row_bitmap <= 16'b0000000000000000;
		15'h3816: char_row_bitmap <= 16'b0000000000000000;
		15'h3817: char_row_bitmap <= 16'b0000000000000000;
		15'h3818: char_row_bitmap <= 16'b0000000000000000;
		15'h3819: char_row_bitmap <= 16'b0000000000000000;
		15'h381a: char_row_bitmap <= 16'b0000000000000000;
		15'h381b: char_row_bitmap <= 16'b0000000000000000;
		15'h381c: char_row_bitmap <= 16'b0000000110000000;
		15'h381d: char_row_bitmap <= 16'b0000000110000000;
		15'h381e: char_row_bitmap <= 16'b0000001111000000;
		15'h381f: char_row_bitmap <= 16'b0000001111000000;
		15'h3820: char_row_bitmap <= 16'b0000011111100000;
		15'h3821: char_row_bitmap <= 16'b0000011111100000;
		15'h3822: char_row_bitmap <= 16'b0000111111110000;
		15'h3823: char_row_bitmap <= 16'b0000111111110000;
		15'h3824: char_row_bitmap <= 16'b0001111111111000;
		15'h3825: char_row_bitmap <= 16'b0001111111111000;
		15'h3826: char_row_bitmap <= 16'b0011111111111100;
		15'h3827: char_row_bitmap <= 16'b0011111111111100;
		15'h3828: char_row_bitmap <= 16'b0111111111111110;
		15'h3829: char_row_bitmap <= 16'b0111111111111110;
		15'h382a: char_row_bitmap <= 16'b1111111111111111;
		15'h382b: char_row_bitmap <= 16'b1111111111111111;
		15'h382c: char_row_bitmap <= 16'b1100000000000000;
		15'h382d: char_row_bitmap <= 16'b1110000000000000;
		15'h382e: char_row_bitmap <= 16'b1111000000000000;
		15'h382f: char_row_bitmap <= 16'b1111100000000000;
		15'h3830: char_row_bitmap <= 16'b1111110000000000;
		15'h3831: char_row_bitmap <= 16'b1111111000000000;
		15'h3832: char_row_bitmap <= 16'b1111111100000000;
		15'h3833: char_row_bitmap <= 16'b1111111110000000;
		15'h3834: char_row_bitmap <= 16'b1111111111000000;
		15'h3835: char_row_bitmap <= 16'b1111111111100000;
		15'h3836: char_row_bitmap <= 16'b1111111111100000;
		15'h3837: char_row_bitmap <= 16'b1111111111000000;
		15'h3838: char_row_bitmap <= 16'b1111111110000000;
		15'h3839: char_row_bitmap <= 16'b1111111100000000;
		15'h383a: char_row_bitmap <= 16'b1111111000000000;
		15'h383b: char_row_bitmap <= 16'b1111110000000000;
		15'h383c: char_row_bitmap <= 16'b1111100000000000;
		15'h383d: char_row_bitmap <= 16'b1111000000000000;
		15'h383e: char_row_bitmap <= 16'b1110000000000000;
		15'h383f: char_row_bitmap <= 16'b1100000000000000;
		15'h3840: char_row_bitmap <= 16'b1111111111111111;
		15'h3841: char_row_bitmap <= 16'b1111111111111111;
		15'h3842: char_row_bitmap <= 16'b1111111111111111;
		15'h3843: char_row_bitmap <= 16'b1111111111111111;
		15'h3844: char_row_bitmap <= 16'b1111111111111111;
		15'h3845: char_row_bitmap <= 16'b1111111111111111;
		15'h3846: char_row_bitmap <= 16'b1111111111111111;
		15'h3847: char_row_bitmap <= 16'b1111111111111111;
		15'h3848: char_row_bitmap <= 16'b1111111111111111;
		15'h3849: char_row_bitmap <= 16'b1111111111111111;
		15'h384a: char_row_bitmap <= 16'b1111111111111111;
		15'h384b: char_row_bitmap <= 16'b1111111111111111;
		15'h384c: char_row_bitmap <= 16'b1111111111111111;
		15'h384d: char_row_bitmap <= 16'b1111111111111111;
		15'h384e: char_row_bitmap <= 16'b1111111111111111;
		15'h384f: char_row_bitmap <= 16'b1111111111111100;
		15'h3850: char_row_bitmap <= 16'b1111111111111000;
		15'h3851: char_row_bitmap <= 16'b1111111111100000;
		15'h3852: char_row_bitmap <= 16'b1111111111000000;
		15'h3853: char_row_bitmap <= 16'b1111111110000000;
		15'h3854: char_row_bitmap <= 16'b1111111111111111;
		15'h3855: char_row_bitmap <= 16'b1111111111111111;
		15'h3856: char_row_bitmap <= 16'b1111111111111111;
		15'h3857: char_row_bitmap <= 16'b1111111111111111;
		15'h3858: char_row_bitmap <= 16'b1111111111111111;
		15'h3859: char_row_bitmap <= 16'b1111111111111111;
		15'h385a: char_row_bitmap <= 16'b1111111111111111;
		15'h385b: char_row_bitmap <= 16'b1111111111111111;
		15'h385c: char_row_bitmap <= 16'b1111111111111111;
		15'h385d: char_row_bitmap <= 16'b1111111111111111;
		15'h385e: char_row_bitmap <= 16'b1111111111111111;
		15'h385f: char_row_bitmap <= 16'b1111111111111111;
		15'h3860: char_row_bitmap <= 16'b1111111111111111;
		15'h3861: char_row_bitmap <= 16'b1111111111111111;
		15'h3862: char_row_bitmap <= 16'b1111111111111100;
		15'h3863: char_row_bitmap <= 16'b1111111111110000;
		15'h3864: char_row_bitmap <= 16'b1111111111000000;
		15'h3865: char_row_bitmap <= 16'b1111111000000000;
		15'h3866: char_row_bitmap <= 16'b1111000000000000;
		15'h3867: char_row_bitmap <= 16'b1100000000000000;
		15'h3868: char_row_bitmap <= 16'b1111111111111111;
		15'h3869: char_row_bitmap <= 16'b1111111111111111;
		15'h386a: char_row_bitmap <= 16'b1111111111111111;
		15'h386b: char_row_bitmap <= 16'b1111111111111111;
		15'h386c: char_row_bitmap <= 16'b1111111111111111;
		15'h386d: char_row_bitmap <= 16'b1111111111111111;
		15'h386e: char_row_bitmap <= 16'b1111111111111111;
		15'h386f: char_row_bitmap <= 16'b1111111111111110;
		15'h3870: char_row_bitmap <= 16'b1111111111111110;
		15'h3871: char_row_bitmap <= 16'b1111111111111100;
		15'h3872: char_row_bitmap <= 16'b1111111111111000;
		15'h3873: char_row_bitmap <= 16'b1111111111111000;
		15'h3874: char_row_bitmap <= 16'b1111111111110000;
		15'h3875: char_row_bitmap <= 16'b1111111111110000;
		15'h3876: char_row_bitmap <= 16'b1111111111100000;
		15'h3877: char_row_bitmap <= 16'b1111111111100000;
		15'h3878: char_row_bitmap <= 16'b1111111111000000;
		15'h3879: char_row_bitmap <= 16'b1111111110000000;
		15'h387a: char_row_bitmap <= 16'b1111111110000000;
		15'h387b: char_row_bitmap <= 16'b1111111100000000;
		15'h387c: char_row_bitmap <= 16'b1111111111111111;
		15'h387d: char_row_bitmap <= 16'b1111111111111100;
		15'h387e: char_row_bitmap <= 16'b1111111111111000;
		15'h387f: char_row_bitmap <= 16'b1111111111110000;
		15'h3880: char_row_bitmap <= 16'b1111111111100000;
		15'h3881: char_row_bitmap <= 16'b1111111111000000;
		15'h3882: char_row_bitmap <= 16'b1111111110000000;
		15'h3883: char_row_bitmap <= 16'b1111111000000000;
		15'h3884: char_row_bitmap <= 16'b1111110000000000;
		15'h3885: char_row_bitmap <= 16'b1111100000000000;
		15'h3886: char_row_bitmap <= 16'b1111000000000000;
		15'h3887: char_row_bitmap <= 16'b1100000000000000;
		15'h3888: char_row_bitmap <= 16'b1000000000000000;
		15'h3889: char_row_bitmap <= 16'b0000000000000000;
		15'h388a: char_row_bitmap <= 16'b0000000000000000;
		15'h388b: char_row_bitmap <= 16'b0000000000000000;
		15'h388c: char_row_bitmap <= 16'b0000000000000000;
		15'h388d: char_row_bitmap <= 16'b0000000000000000;
		15'h388e: char_row_bitmap <= 16'b0000000000000000;
		15'h388f: char_row_bitmap <= 16'b0000000000000000;
		15'h3890: char_row_bitmap <= 16'b1111111111111111;
		15'h3891: char_row_bitmap <= 16'b1111111111111110;
		15'h3892: char_row_bitmap <= 16'b1111111111111110;
		15'h3893: char_row_bitmap <= 16'b1111111111111110;
		15'h3894: char_row_bitmap <= 16'b1111111111111100;
		15'h3895: char_row_bitmap <= 16'b1111111111111100;
		15'h3896: char_row_bitmap <= 16'b1111111111111000;
		15'h3897: char_row_bitmap <= 16'b1111111111111000;
		15'h3898: char_row_bitmap <= 16'b1111111111111000;
		15'h3899: char_row_bitmap <= 16'b1111111111110000;
		15'h389a: char_row_bitmap <= 16'b1111111111110000;
		15'h389b: char_row_bitmap <= 16'b1111111111100000;
		15'h389c: char_row_bitmap <= 16'b1111111111100000;
		15'h389d: char_row_bitmap <= 16'b1111111111100000;
		15'h389e: char_row_bitmap <= 16'b1111111111000000;
		15'h389f: char_row_bitmap <= 16'b1111111111000000;
		15'h38a0: char_row_bitmap <= 16'b1111111110000000;
		15'h38a1: char_row_bitmap <= 16'b1111111110000000;
		15'h38a2: char_row_bitmap <= 16'b1111111110000000;
		15'h38a3: char_row_bitmap <= 16'b1111111100000000;
		15'h38a4: char_row_bitmap <= 16'b1111111111111111;
		15'h38a5: char_row_bitmap <= 16'b1111111111111110;
		15'h38a6: char_row_bitmap <= 16'b1111111111111100;
		15'h38a7: char_row_bitmap <= 16'b1111111111111000;
		15'h38a8: char_row_bitmap <= 16'b1111111111110000;
		15'h38a9: char_row_bitmap <= 16'b1111111111110000;
		15'h38aa: char_row_bitmap <= 16'b1111111111100000;
		15'h38ab: char_row_bitmap <= 16'b1111111111000000;
		15'h38ac: char_row_bitmap <= 16'b1111111110000000;
		15'h38ad: char_row_bitmap <= 16'b1111111100000000;
		15'h38ae: char_row_bitmap <= 16'b1111111100000000;
		15'h38af: char_row_bitmap <= 16'b1111111000000000;
		15'h38b0: char_row_bitmap <= 16'b1111110000000000;
		15'h38b1: char_row_bitmap <= 16'b1111100000000000;
		15'h38b2: char_row_bitmap <= 16'b1111000000000000;
		15'h38b3: char_row_bitmap <= 16'b1111000000000000;
		15'h38b4: char_row_bitmap <= 16'b1110000000000000;
		15'h38b5: char_row_bitmap <= 16'b1100000000000000;
		15'h38b6: char_row_bitmap <= 16'b1100000000000000;
		15'h38b7: char_row_bitmap <= 16'b1000000000000000;
		15'h38b8: char_row_bitmap <= 16'b0000000011111111;
		15'h38b9: char_row_bitmap <= 16'b0000000000111111;
		15'h38ba: char_row_bitmap <= 16'b0000000000011111;
		15'h38bb: char_row_bitmap <= 16'b0000000000000111;
		15'h38bc: char_row_bitmap <= 16'b0000000000000011;
		15'h38bd: char_row_bitmap <= 16'b0000000000000001;
		15'h38be: char_row_bitmap <= 16'b0000000000000000;
		15'h38bf: char_row_bitmap <= 16'b0000000000000000;
		15'h38c0: char_row_bitmap <= 16'b0000000000000000;
		15'h38c1: char_row_bitmap <= 16'b0000000000000000;
		15'h38c2: char_row_bitmap <= 16'b0000000000000000;
		15'h38c3: char_row_bitmap <= 16'b0000000000000000;
		15'h38c4: char_row_bitmap <= 16'b0000000000000000;
		15'h38c5: char_row_bitmap <= 16'b0000000000000000;
		15'h38c6: char_row_bitmap <= 16'b0000000000000000;
		15'h38c7: char_row_bitmap <= 16'b0000000000000000;
		15'h38c8: char_row_bitmap <= 16'b0000000000000000;
		15'h38c9: char_row_bitmap <= 16'b0000000000000000;
		15'h38ca: char_row_bitmap <= 16'b0000000000000000;
		15'h38cb: char_row_bitmap <= 16'b0000000000000000;
		15'h38cc: char_row_bitmap <= 16'b0111111111111111;
		15'h38cd: char_row_bitmap <= 16'b0001111111111111;
		15'h38ce: char_row_bitmap <= 16'b0000001111111111;
		15'h38cf: char_row_bitmap <= 16'b0000000001111111;
		15'h38d0: char_row_bitmap <= 16'b0000000000001111;
		15'h38d1: char_row_bitmap <= 16'b0000000000000011;
		15'h38d2: char_row_bitmap <= 16'b0000000000000000;
		15'h38d3: char_row_bitmap <= 16'b0000000000000000;
		15'h38d4: char_row_bitmap <= 16'b0000000000000000;
		15'h38d5: char_row_bitmap <= 16'b0000000000000000;
		15'h38d6: char_row_bitmap <= 16'b0000000000000000;
		15'h38d7: char_row_bitmap <= 16'b0000000000000000;
		15'h38d8: char_row_bitmap <= 16'b0000000000000000;
		15'h38d9: char_row_bitmap <= 16'b0000000000000000;
		15'h38da: char_row_bitmap <= 16'b0000000000000000;
		15'h38db: char_row_bitmap <= 16'b0000000000000000;
		15'h38dc: char_row_bitmap <= 16'b0000000000000000;
		15'h38dd: char_row_bitmap <= 16'b0000000000000000;
		15'h38de: char_row_bitmap <= 16'b0000000000000000;
		15'h38df: char_row_bitmap <= 16'b0000000000000000;
		15'h38e0: char_row_bitmap <= 16'b0000000011111111;
		15'h38e1: char_row_bitmap <= 16'b0000000001111111;
		15'h38e2: char_row_bitmap <= 16'b0000000001111111;
		15'h38e3: char_row_bitmap <= 16'b0000000000111111;
		15'h38e4: char_row_bitmap <= 16'b0000000000011111;
		15'h38e5: char_row_bitmap <= 16'b0000000000011111;
		15'h38e6: char_row_bitmap <= 16'b0000000000001111;
		15'h38e7: char_row_bitmap <= 16'b0000000000001111;
		15'h38e8: char_row_bitmap <= 16'b0000000000000111;
		15'h38e9: char_row_bitmap <= 16'b0000000000000111;
		15'h38ea: char_row_bitmap <= 16'b0000000000000011;
		15'h38eb: char_row_bitmap <= 16'b0000000000000011;
		15'h38ec: char_row_bitmap <= 16'b0000000000000001;
		15'h38ed: char_row_bitmap <= 16'b0000000000000001;
		15'h38ee: char_row_bitmap <= 16'b0000000000000000;
		15'h38ef: char_row_bitmap <= 16'b0000000000000000;
		15'h38f0: char_row_bitmap <= 16'b0000000000000000;
		15'h38f1: char_row_bitmap <= 16'b0000000000000000;
		15'h38f2: char_row_bitmap <= 16'b0000000000000000;
		15'h38f3: char_row_bitmap <= 16'b0000000000000000;
		15'h38f4: char_row_bitmap <= 16'b0111111111111111;
		15'h38f5: char_row_bitmap <= 16'b0011111111111111;
		15'h38f6: char_row_bitmap <= 16'b0001111111111111;
		15'h38f7: char_row_bitmap <= 16'b0000111111111111;
		15'h38f8: char_row_bitmap <= 16'b0000011111111111;
		15'h38f9: char_row_bitmap <= 16'b0000001111111111;
		15'h38fa: char_row_bitmap <= 16'b0000000111111111;
		15'h38fb: char_row_bitmap <= 16'b0000000001111111;
		15'h38fc: char_row_bitmap <= 16'b0000000000111111;
		15'h38fd: char_row_bitmap <= 16'b0000000000011111;
		15'h38fe: char_row_bitmap <= 16'b0000000000001111;
		15'h38ff: char_row_bitmap <= 16'b0000000000000011;
		15'h3900: char_row_bitmap <= 16'b0000000000000001;
		15'h3901: char_row_bitmap <= 16'b0000000000000000;
		15'h3902: char_row_bitmap <= 16'b0000000000000000;
		15'h3903: char_row_bitmap <= 16'b0000000000000000;
		15'h3904: char_row_bitmap <= 16'b0000000000000000;
		15'h3905: char_row_bitmap <= 16'b0000000000000000;
		15'h3906: char_row_bitmap <= 16'b0000000000000000;
		15'h3907: char_row_bitmap <= 16'b0000000000000000;
		15'h3908: char_row_bitmap <= 16'b0000000011111111;
		15'h3909: char_row_bitmap <= 16'b0000000001111111;
		15'h390a: char_row_bitmap <= 16'b0000000001111111;
		15'h390b: char_row_bitmap <= 16'b0000000001111111;
		15'h390c: char_row_bitmap <= 16'b0000000000111111;
		15'h390d: char_row_bitmap <= 16'b0000000000111111;
		15'h390e: char_row_bitmap <= 16'b0000000000011111;
		15'h390f: char_row_bitmap <= 16'b0000000000011111;
		15'h3910: char_row_bitmap <= 16'b0000000000011111;
		15'h3911: char_row_bitmap <= 16'b0000000000001111;
		15'h3912: char_row_bitmap <= 16'b0000000000001111;
		15'h3913: char_row_bitmap <= 16'b0000000000001111;
		15'h3914: char_row_bitmap <= 16'b0000000000000111;
		15'h3915: char_row_bitmap <= 16'b0000000000000111;
		15'h3916: char_row_bitmap <= 16'b0000000000000111;
		15'h3917: char_row_bitmap <= 16'b0000000000000011;
		15'h3918: char_row_bitmap <= 16'b0000000000000011;
		15'h3919: char_row_bitmap <= 16'b0000000000000011;
		15'h391a: char_row_bitmap <= 16'b0000000000000001;
		15'h391b: char_row_bitmap <= 16'b0000000000000001;
		15'h391c: char_row_bitmap <= 16'b1111111111111111;
		15'h391d: char_row_bitmap <= 16'b1111111111111111;
		15'h391e: char_row_bitmap <= 16'b1111111111111111;
		15'h391f: char_row_bitmap <= 16'b1111111111111111;
		15'h3920: char_row_bitmap <= 16'b1111111111111111;
		15'h3921: char_row_bitmap <= 16'b1111111111111111;
		15'h3922: char_row_bitmap <= 16'b0111111111111111;
		15'h3923: char_row_bitmap <= 16'b0001111111111111;
		15'h3924: char_row_bitmap <= 16'b0000011111111111;
		15'h3925: char_row_bitmap <= 16'b0000000111111111;
		15'h3926: char_row_bitmap <= 16'b0000000001111111;
		15'h3927: char_row_bitmap <= 16'b0000000000011111;
		15'h3928: char_row_bitmap <= 16'b0000000000000111;
		15'h3929: char_row_bitmap <= 16'b0000000000000001;
		15'h392a: char_row_bitmap <= 16'b0000000000000000;
		15'h392b: char_row_bitmap <= 16'b0000000000000000;
		15'h392c: char_row_bitmap <= 16'b0000000000000000;
		15'h392d: char_row_bitmap <= 16'b0000000000000000;
		15'h392e: char_row_bitmap <= 16'b0000000000000000;
		15'h392f: char_row_bitmap <= 16'b0000000000000000;
		15'h3930: char_row_bitmap <= 16'b0000000000000000;
		15'h3931: char_row_bitmap <= 16'b0000000000000001;
		15'h3932: char_row_bitmap <= 16'b0000000000000011;
		15'h3933: char_row_bitmap <= 16'b0000000000000111;
		15'h3934: char_row_bitmap <= 16'b0000000000001111;
		15'h3935: char_row_bitmap <= 16'b0000000000011111;
		15'h3936: char_row_bitmap <= 16'b0000000000111111;
		15'h3937: char_row_bitmap <= 16'b0000000001111111;
		15'h3938: char_row_bitmap <= 16'b0000000011111111;
		15'h3939: char_row_bitmap <= 16'b0000000111111111;
		15'h393a: char_row_bitmap <= 16'b0000000111111111;
		15'h393b: char_row_bitmap <= 16'b0000000011111111;
		15'h393c: char_row_bitmap <= 16'b0000000001111111;
		15'h393d: char_row_bitmap <= 16'b0000000000111111;
		15'h393e: char_row_bitmap <= 16'b0000000000011111;
		15'h393f: char_row_bitmap <= 16'b0000000000001111;
		15'h3940: char_row_bitmap <= 16'b0000000000000111;
		15'h3941: char_row_bitmap <= 16'b0000000000000011;
		15'h3942: char_row_bitmap <= 16'b0000000000000001;
		15'h3943: char_row_bitmap <= 16'b0000000000000000;
		15'h3944: char_row_bitmap <= 16'b0000000000000000;
		15'h3945: char_row_bitmap <= 16'b0000000000000000;
		15'h3946: char_row_bitmap <= 16'b0000000000000000;
		15'h3947: char_row_bitmap <= 16'b0000000000000000;
		15'h3948: char_row_bitmap <= 16'b0000000000000000;
		15'h3949: char_row_bitmap <= 16'b0000000000000000;
		15'h394a: char_row_bitmap <= 16'b0000000000000000;
		15'h394b: char_row_bitmap <= 16'b0000000000000000;
		15'h394c: char_row_bitmap <= 16'b0000000000000000;
		15'h394d: char_row_bitmap <= 16'b0000000000000000;
		15'h394e: char_row_bitmap <= 16'b0000000000000000;
		15'h394f: char_row_bitmap <= 16'b0000000000000000;
		15'h3950: char_row_bitmap <= 16'b0000000000000000;
		15'h3951: char_row_bitmap <= 16'b0000000110000000;
		15'h3952: char_row_bitmap <= 16'b0000001111000000;
		15'h3953: char_row_bitmap <= 16'b0000011111100000;
		15'h3954: char_row_bitmap <= 16'b0000111111110000;
		15'h3955: char_row_bitmap <= 16'b0001111111111000;
		15'h3956: char_row_bitmap <= 16'b0011111111111100;
		15'h3957: char_row_bitmap <= 16'b0111111111111110;
		15'h3958: char_row_bitmap <= 16'b1111111111111111;
		15'h3959: char_row_bitmap <= 16'b1111111111111111;
		15'h395a: char_row_bitmap <= 16'b0111111111111110;
		15'h395b: char_row_bitmap <= 16'b0111111111111110;
		15'h395c: char_row_bitmap <= 16'b0011111111111100;
		15'h395d: char_row_bitmap <= 16'b0011111111111100;
		15'h395e: char_row_bitmap <= 16'b0001111111111000;
		15'h395f: char_row_bitmap <= 16'b0001111111111000;
		15'h3960: char_row_bitmap <= 16'b0000111111110000;
		15'h3961: char_row_bitmap <= 16'b0000111111110000;
		15'h3962: char_row_bitmap <= 16'b0000011111100000;
		15'h3963: char_row_bitmap <= 16'b0000011111100000;
		15'h3964: char_row_bitmap <= 16'b0000001111000000;
		15'h3965: char_row_bitmap <= 16'b0000001111000000;
		15'h3966: char_row_bitmap <= 16'b0000000110000000;
		15'h3967: char_row_bitmap <= 16'b0000000110000000;
		15'h3968: char_row_bitmap <= 16'b0000000000000000;
		15'h3969: char_row_bitmap <= 16'b0000000000000000;
		15'h396a: char_row_bitmap <= 16'b0000000000000000;
		15'h396b: char_row_bitmap <= 16'b0000000000000000;
		15'h396c: char_row_bitmap <= 16'b0000000000000011;
		15'h396d: char_row_bitmap <= 16'b0000000000000111;
		15'h396e: char_row_bitmap <= 16'b0000000000001111;
		15'h396f: char_row_bitmap <= 16'b0000000000011111;
		15'h3970: char_row_bitmap <= 16'b0000000000111111;
		15'h3971: char_row_bitmap <= 16'b0000000001111111;
		15'h3972: char_row_bitmap <= 16'b0000000011111111;
		15'h3973: char_row_bitmap <= 16'b0000000111111111;
		15'h3974: char_row_bitmap <= 16'b0000001111111111;
		15'h3975: char_row_bitmap <= 16'b0000011111111111;
		15'h3976: char_row_bitmap <= 16'b0000011111111111;
		15'h3977: char_row_bitmap <= 16'b0000001111111111;
		15'h3978: char_row_bitmap <= 16'b0000000111111111;
		15'h3979: char_row_bitmap <= 16'b0000000011111111;
		15'h397a: char_row_bitmap <= 16'b0000000001111111;
		15'h397b: char_row_bitmap <= 16'b0000000000111111;
		15'h397c: char_row_bitmap <= 16'b0000000000011111;
		15'h397d: char_row_bitmap <= 16'b0000000000001111;
		15'h397e: char_row_bitmap <= 16'b0000000000000111;
		15'h397f: char_row_bitmap <= 16'b0000000000000011;
		15'h3980: char_row_bitmap <= 16'b1100000000000000;
		15'h3981: char_row_bitmap <= 16'b1100000000000000;
		15'h3982: char_row_bitmap <= 16'b1100000000000000;
		15'h3983: char_row_bitmap <= 16'b1100000000000000;
		15'h3984: char_row_bitmap <= 16'b1100000000000000;
		15'h3985: char_row_bitmap <= 16'b1100000000000000;
		15'h3986: char_row_bitmap <= 16'b1100000000000000;
		15'h3987: char_row_bitmap <= 16'b1100000000000000;
		15'h3988: char_row_bitmap <= 16'b1100000000000000;
		15'h3989: char_row_bitmap <= 16'b1100000000000000;
		15'h398a: char_row_bitmap <= 16'b1100000000000000;
		15'h398b: char_row_bitmap <= 16'b1100000000000000;
		15'h398c: char_row_bitmap <= 16'b1100000000000000;
		15'h398d: char_row_bitmap <= 16'b1100000000000000;
		15'h398e: char_row_bitmap <= 16'b1100000000000000;
		15'h398f: char_row_bitmap <= 16'b1100000000000000;
		15'h3990: char_row_bitmap <= 16'b1100000000000000;
		15'h3991: char_row_bitmap <= 16'b1100000000000000;
		15'h3992: char_row_bitmap <= 16'b1100000000000000;
		15'h3993: char_row_bitmap <= 16'b1100000000000000;
		15'h3994: char_row_bitmap <= 16'b1111000000000000;
		15'h3995: char_row_bitmap <= 16'b1111000000000000;
		15'h3996: char_row_bitmap <= 16'b1111000000000000;
		15'h3997: char_row_bitmap <= 16'b1111000000000000;
		15'h3998: char_row_bitmap <= 16'b1111000000000000;
		15'h3999: char_row_bitmap <= 16'b1111000000000000;
		15'h399a: char_row_bitmap <= 16'b1111000000000000;
		15'h399b: char_row_bitmap <= 16'b1111000000000000;
		15'h399c: char_row_bitmap <= 16'b1111000000000000;
		15'h399d: char_row_bitmap <= 16'b1111000000000000;
		15'h399e: char_row_bitmap <= 16'b1111000000000000;
		15'h399f: char_row_bitmap <= 16'b1111000000000000;
		15'h39a0: char_row_bitmap <= 16'b1111000000000000;
		15'h39a1: char_row_bitmap <= 16'b1111000000000000;
		15'h39a2: char_row_bitmap <= 16'b1111000000000000;
		15'h39a3: char_row_bitmap <= 16'b1111000000000000;
		15'h39a4: char_row_bitmap <= 16'b1111000000000000;
		15'h39a5: char_row_bitmap <= 16'b1111000000000000;
		15'h39a6: char_row_bitmap <= 16'b1111000000000000;
		15'h39a7: char_row_bitmap <= 16'b1111000000000000;
		15'h39a8: char_row_bitmap <= 16'b1111110000000000;
		15'h39a9: char_row_bitmap <= 16'b1111110000000000;
		15'h39aa: char_row_bitmap <= 16'b1111110000000000;
		15'h39ab: char_row_bitmap <= 16'b1111110000000000;
		15'h39ac: char_row_bitmap <= 16'b1111110000000000;
		15'h39ad: char_row_bitmap <= 16'b1111110000000000;
		15'h39ae: char_row_bitmap <= 16'b1111110000000000;
		15'h39af: char_row_bitmap <= 16'b1111110000000000;
		15'h39b0: char_row_bitmap <= 16'b1111110000000000;
		15'h39b1: char_row_bitmap <= 16'b1111110000000000;
		15'h39b2: char_row_bitmap <= 16'b1111110000000000;
		15'h39b3: char_row_bitmap <= 16'b1111110000000000;
		15'h39b4: char_row_bitmap <= 16'b1111110000000000;
		15'h39b5: char_row_bitmap <= 16'b1111110000000000;
		15'h39b6: char_row_bitmap <= 16'b1111110000000000;
		15'h39b7: char_row_bitmap <= 16'b1111110000000000;
		15'h39b8: char_row_bitmap <= 16'b1111110000000000;
		15'h39b9: char_row_bitmap <= 16'b1111110000000000;
		15'h39ba: char_row_bitmap <= 16'b1111110000000000;
		15'h39bb: char_row_bitmap <= 16'b1111110000000000;
		15'h39bc: char_row_bitmap <= 16'b1111111100000000;
		15'h39bd: char_row_bitmap <= 16'b1111111100000000;
		15'h39be: char_row_bitmap <= 16'b1111111100000000;
		15'h39bf: char_row_bitmap <= 16'b1111111100000000;
		15'h39c0: char_row_bitmap <= 16'b1111111100000000;
		15'h39c1: char_row_bitmap <= 16'b1111111100000000;
		15'h39c2: char_row_bitmap <= 16'b1111111100000000;
		15'h39c3: char_row_bitmap <= 16'b1111111100000000;
		15'h39c4: char_row_bitmap <= 16'b1111111100000000;
		15'h39c5: char_row_bitmap <= 16'b1111111100000000;
		15'h39c6: char_row_bitmap <= 16'b1111111100000000;
		15'h39c7: char_row_bitmap <= 16'b1111111100000000;
		15'h39c8: char_row_bitmap <= 16'b1111111100000000;
		15'h39c9: char_row_bitmap <= 16'b1111111100000000;
		15'h39ca: char_row_bitmap <= 16'b1111111100000000;
		15'h39cb: char_row_bitmap <= 16'b1111111100000000;
		15'h39cc: char_row_bitmap <= 16'b1111111100000000;
		15'h39cd: char_row_bitmap <= 16'b1111111100000000;
		15'h39ce: char_row_bitmap <= 16'b1111111100000000;
		15'h39cf: char_row_bitmap <= 16'b1111111100000000;
		15'h39d0: char_row_bitmap <= 16'b1111111111000000;
		15'h39d1: char_row_bitmap <= 16'b1111111111000000;
		15'h39d2: char_row_bitmap <= 16'b1111111111000000;
		15'h39d3: char_row_bitmap <= 16'b1111111111000000;
		15'h39d4: char_row_bitmap <= 16'b1111111111000000;
		15'h39d5: char_row_bitmap <= 16'b1111111111000000;
		15'h39d6: char_row_bitmap <= 16'b1111111111000000;
		15'h39d7: char_row_bitmap <= 16'b1111111111000000;
		15'h39d8: char_row_bitmap <= 16'b1111111111000000;
		15'h39d9: char_row_bitmap <= 16'b1111111111000000;
		15'h39da: char_row_bitmap <= 16'b1111111111000000;
		15'h39db: char_row_bitmap <= 16'b1111111111000000;
		15'h39dc: char_row_bitmap <= 16'b1111111111000000;
		15'h39dd: char_row_bitmap <= 16'b1111111111000000;
		15'h39de: char_row_bitmap <= 16'b1111111111000000;
		15'h39df: char_row_bitmap <= 16'b1111111111000000;
		15'h39e0: char_row_bitmap <= 16'b1111111111000000;
		15'h39e1: char_row_bitmap <= 16'b1111111111000000;
		15'h39e2: char_row_bitmap <= 16'b1111111111000000;
		15'h39e3: char_row_bitmap <= 16'b1111111111000000;
		15'h39e4: char_row_bitmap <= 16'b1111111111110000;
		15'h39e5: char_row_bitmap <= 16'b1111111111110000;
		15'h39e6: char_row_bitmap <= 16'b1111111111110000;
		15'h39e7: char_row_bitmap <= 16'b1111111111110000;
		15'h39e8: char_row_bitmap <= 16'b1111111111110000;
		15'h39e9: char_row_bitmap <= 16'b1111111111110000;
		15'h39ea: char_row_bitmap <= 16'b1111111111110000;
		15'h39eb: char_row_bitmap <= 16'b1111111111110000;
		15'h39ec: char_row_bitmap <= 16'b1111111111110000;
		15'h39ed: char_row_bitmap <= 16'b1111111111110000;
		15'h39ee: char_row_bitmap <= 16'b1111111111110000;
		15'h39ef: char_row_bitmap <= 16'b1111111111110000;
		15'h39f0: char_row_bitmap <= 16'b1111111111110000;
		15'h39f1: char_row_bitmap <= 16'b1111111111110000;
		15'h39f2: char_row_bitmap <= 16'b1111111111110000;
		15'h39f3: char_row_bitmap <= 16'b1111111111110000;
		15'h39f4: char_row_bitmap <= 16'b1111111111110000;
		15'h39f5: char_row_bitmap <= 16'b1111111111110000;
		15'h39f6: char_row_bitmap <= 16'b1111111111110000;
		15'h39f7: char_row_bitmap <= 16'b1111111111110000;
		15'h39f8: char_row_bitmap <= 16'b1111111111111100;
		15'h39f9: char_row_bitmap <= 16'b1111111111111100;
		15'h39fa: char_row_bitmap <= 16'b1111111111111100;
		15'h39fb: char_row_bitmap <= 16'b1111111111111100;
		15'h39fc: char_row_bitmap <= 16'b1111111111111100;
		15'h39fd: char_row_bitmap <= 16'b1111111111111100;
		15'h39fe: char_row_bitmap <= 16'b1111111111111100;
		15'h39ff: char_row_bitmap <= 16'b1111111111111100;
		15'h3a00: char_row_bitmap <= 16'b1111111111111100;
		15'h3a01: char_row_bitmap <= 16'b1111111111111100;
		15'h3a02: char_row_bitmap <= 16'b1111111111111100;
		15'h3a03: char_row_bitmap <= 16'b1111111111111100;
		15'h3a04: char_row_bitmap <= 16'b1111111111111100;
		15'h3a05: char_row_bitmap <= 16'b1111111111111100;
		15'h3a06: char_row_bitmap <= 16'b1111111111111100;
		15'h3a07: char_row_bitmap <= 16'b1111111111111100;
		15'h3a08: char_row_bitmap <= 16'b1111111111111100;
		15'h3a09: char_row_bitmap <= 16'b1111111111111100;
		15'h3a0a: char_row_bitmap <= 16'b1111111111111100;
		15'h3a0b: char_row_bitmap <= 16'b1111111111111100;
		15'h3a0c: char_row_bitmap <= 16'b1111111111111111;
		15'h3a0d: char_row_bitmap <= 16'b1111111111111111;
		15'h3a0e: char_row_bitmap <= 16'b1111111111111111;
		15'h3a0f: char_row_bitmap <= 16'b1111111111111111;
		15'h3a10: char_row_bitmap <= 16'b1111111111111111;
		15'h3a11: char_row_bitmap <= 16'b1111111111111111;
		15'h3a12: char_row_bitmap <= 16'b1111111111111111;
		15'h3a13: char_row_bitmap <= 16'b1111111111111111;
		15'h3a14: char_row_bitmap <= 16'b1111111111111111;
		15'h3a15: char_row_bitmap <= 16'b1111111111111111;
		15'h3a16: char_row_bitmap <= 16'b1111111111111111;
		15'h3a17: char_row_bitmap <= 16'b1111111111111111;
		15'h3a18: char_row_bitmap <= 16'b1111111111111111;
		15'h3a19: char_row_bitmap <= 16'b1111111111111111;
		15'h3a1a: char_row_bitmap <= 16'b1111111111111111;
		15'h3a1b: char_row_bitmap <= 16'b1111111111111111;
		15'h3a1c: char_row_bitmap <= 16'b1111111111111111;
		15'h3a1d: char_row_bitmap <= 16'b1111111111111111;
		15'h3a1e: char_row_bitmap <= 16'b1111111111111111;
		15'h3a1f: char_row_bitmap <= 16'b1111111111111111;
		15'h3a20: char_row_bitmap <= 16'b1000000000000000;
		15'h3a21: char_row_bitmap <= 16'b1000000000000000;
		15'h3a22: char_row_bitmap <= 16'b1000000000000000;
		15'h3a23: char_row_bitmap <= 16'b1000000000000000;
		15'h3a24: char_row_bitmap <= 16'b1000000000000000;
		15'h3a25: char_row_bitmap <= 16'b1000000000000000;
		15'h3a26: char_row_bitmap <= 16'b1000000000000000;
		15'h3a27: char_row_bitmap <= 16'b1000000000000000;
		15'h3a28: char_row_bitmap <= 16'b1000000000000000;
		15'h3a29: char_row_bitmap <= 16'b1000000000000000;
		15'h3a2a: char_row_bitmap <= 16'b1000000000000000;
		15'h3a2b: char_row_bitmap <= 16'b1000000000000000;
		15'h3a2c: char_row_bitmap <= 16'b1000000000000000;
		15'h3a2d: char_row_bitmap <= 16'b1000000000000000;
		15'h3a2e: char_row_bitmap <= 16'b1000000000000000;
		15'h3a2f: char_row_bitmap <= 16'b1000000000000000;
		15'h3a30: char_row_bitmap <= 16'b1000000000000000;
		15'h3a31: char_row_bitmap <= 16'b1000000000000000;
		15'h3a32: char_row_bitmap <= 16'b0000000000000000;
		15'h3a33: char_row_bitmap <= 16'b0000000000000000;
		15'h3a34: char_row_bitmap <= 16'b1111000000000000;
		15'h3a35: char_row_bitmap <= 16'b1111000000000000;
		15'h3a36: char_row_bitmap <= 16'b1111000000000000;
		15'h3a37: char_row_bitmap <= 16'b1111000000000000;
		15'h3a38: char_row_bitmap <= 16'b1111000000000000;
		15'h3a39: char_row_bitmap <= 16'b1111000000000000;
		15'h3a3a: char_row_bitmap <= 16'b1111000000000000;
		15'h3a3b: char_row_bitmap <= 16'b1111000000000000;
		15'h3a3c: char_row_bitmap <= 16'b1111000000000000;
		15'h3a3d: char_row_bitmap <= 16'b1111000000000000;
		15'h3a3e: char_row_bitmap <= 16'b1111000000000000;
		15'h3a3f: char_row_bitmap <= 16'b1111000000000000;
		15'h3a40: char_row_bitmap <= 16'b1111000000000000;
		15'h3a41: char_row_bitmap <= 16'b1111000000000000;
		15'h3a42: char_row_bitmap <= 16'b1111000000000000;
		15'h3a43: char_row_bitmap <= 16'b1111000000000000;
		15'h3a44: char_row_bitmap <= 16'b1111000000000000;
		15'h3a45: char_row_bitmap <= 16'b1111000000000000;
		15'h3a46: char_row_bitmap <= 16'b0000000000000000;
		15'h3a47: char_row_bitmap <= 16'b0000000000000000;
		15'h3a48: char_row_bitmap <= 16'b1111110000000000;
		15'h3a49: char_row_bitmap <= 16'b1111110000000000;
		15'h3a4a: char_row_bitmap <= 16'b1111110000000000;
		15'h3a4b: char_row_bitmap <= 16'b1111110000000000;
		15'h3a4c: char_row_bitmap <= 16'b1111110000000000;
		15'h3a4d: char_row_bitmap <= 16'b1111110000000000;
		15'h3a4e: char_row_bitmap <= 16'b1111110000000000;
		15'h3a4f: char_row_bitmap <= 16'b1111110000000000;
		15'h3a50: char_row_bitmap <= 16'b1111110000000000;
		15'h3a51: char_row_bitmap <= 16'b1111110000000000;
		15'h3a52: char_row_bitmap <= 16'b1111110000000000;
		15'h3a53: char_row_bitmap <= 16'b1111110000000000;
		15'h3a54: char_row_bitmap <= 16'b1111110000000000;
		15'h3a55: char_row_bitmap <= 16'b1111110000000000;
		15'h3a56: char_row_bitmap <= 16'b1111110000000000;
		15'h3a57: char_row_bitmap <= 16'b1111110000000000;
		15'h3a58: char_row_bitmap <= 16'b1111110000000000;
		15'h3a59: char_row_bitmap <= 16'b1111110000000000;
		15'h3a5a: char_row_bitmap <= 16'b0000000000000000;
		15'h3a5b: char_row_bitmap <= 16'b0000000000000000;
		15'h3a5c: char_row_bitmap <= 16'b1111111100000000;
		15'h3a5d: char_row_bitmap <= 16'b1111111100000000;
		15'h3a5e: char_row_bitmap <= 16'b1111111100000000;
		15'h3a5f: char_row_bitmap <= 16'b1111111100000000;
		15'h3a60: char_row_bitmap <= 16'b1111111100000000;
		15'h3a61: char_row_bitmap <= 16'b1111111100000000;
		15'h3a62: char_row_bitmap <= 16'b1111111100000000;
		15'h3a63: char_row_bitmap <= 16'b1111111100000000;
		15'h3a64: char_row_bitmap <= 16'b1111111100000000;
		15'h3a65: char_row_bitmap <= 16'b1111111100000000;
		15'h3a66: char_row_bitmap <= 16'b1111111100000000;
		15'h3a67: char_row_bitmap <= 16'b1111111100000000;
		15'h3a68: char_row_bitmap <= 16'b1111111100000000;
		15'h3a69: char_row_bitmap <= 16'b1111111100000000;
		15'h3a6a: char_row_bitmap <= 16'b1111111100000000;
		15'h3a6b: char_row_bitmap <= 16'b1111111100000000;
		15'h3a6c: char_row_bitmap <= 16'b1111111100000000;
		15'h3a6d: char_row_bitmap <= 16'b1111111100000000;
		15'h3a6e: char_row_bitmap <= 16'b0000000000000000;
		15'h3a6f: char_row_bitmap <= 16'b0000000000000000;
		15'h3a70: char_row_bitmap <= 16'b1111111111000000;
		15'h3a71: char_row_bitmap <= 16'b1111111111000000;
		15'h3a72: char_row_bitmap <= 16'b1111111111000000;
		15'h3a73: char_row_bitmap <= 16'b1111111111000000;
		15'h3a74: char_row_bitmap <= 16'b1111111111000000;
		15'h3a75: char_row_bitmap <= 16'b1111111111000000;
		15'h3a76: char_row_bitmap <= 16'b1111111111000000;
		15'h3a77: char_row_bitmap <= 16'b1111111111000000;
		15'h3a78: char_row_bitmap <= 16'b1111111111000000;
		15'h3a79: char_row_bitmap <= 16'b1111111111000000;
		15'h3a7a: char_row_bitmap <= 16'b1111111111000000;
		15'h3a7b: char_row_bitmap <= 16'b1111111111000000;
		15'h3a7c: char_row_bitmap <= 16'b1111111111000000;
		15'h3a7d: char_row_bitmap <= 16'b1111111111000000;
		15'h3a7e: char_row_bitmap <= 16'b1111111111000000;
		15'h3a7f: char_row_bitmap <= 16'b1111111111000000;
		15'h3a80: char_row_bitmap <= 16'b1111111111000000;
		15'h3a81: char_row_bitmap <= 16'b1111111111000000;
		15'h3a82: char_row_bitmap <= 16'b0000000000000000;
		15'h3a83: char_row_bitmap <= 16'b0000000000000000;
		15'h3a84: char_row_bitmap <= 16'b1111111111110000;
		15'h3a85: char_row_bitmap <= 16'b1111111111110000;
		15'h3a86: char_row_bitmap <= 16'b1111111111110000;
		15'h3a87: char_row_bitmap <= 16'b1111111111110000;
		15'h3a88: char_row_bitmap <= 16'b1111111111110000;
		15'h3a89: char_row_bitmap <= 16'b1111111111110000;
		15'h3a8a: char_row_bitmap <= 16'b1111111111110000;
		15'h3a8b: char_row_bitmap <= 16'b1111111111110000;
		15'h3a8c: char_row_bitmap <= 16'b1111111111110000;
		15'h3a8d: char_row_bitmap <= 16'b1111111111110000;
		15'h3a8e: char_row_bitmap <= 16'b1111111111110000;
		15'h3a8f: char_row_bitmap <= 16'b1111111111110000;
		15'h3a90: char_row_bitmap <= 16'b1111111111110000;
		15'h3a91: char_row_bitmap <= 16'b1111111111110000;
		15'h3a92: char_row_bitmap <= 16'b1111111111110000;
		15'h3a93: char_row_bitmap <= 16'b1111111111110000;
		15'h3a94: char_row_bitmap <= 16'b1111111111110000;
		15'h3a95: char_row_bitmap <= 16'b1111111111110000;
		15'h3a96: char_row_bitmap <= 16'b0000000000000000;
		15'h3a97: char_row_bitmap <= 16'b0000000000000000;
		15'h3a98: char_row_bitmap <= 16'b1111111111111100;
		15'h3a99: char_row_bitmap <= 16'b1111111111111100;
		15'h3a9a: char_row_bitmap <= 16'b1111111111111100;
		15'h3a9b: char_row_bitmap <= 16'b1111111111111100;
		15'h3a9c: char_row_bitmap <= 16'b1111111111111100;
		15'h3a9d: char_row_bitmap <= 16'b1111111111111100;
		15'h3a9e: char_row_bitmap <= 16'b1111111111111100;
		15'h3a9f: char_row_bitmap <= 16'b1111111111111100;
		15'h3aa0: char_row_bitmap <= 16'b1111111111111100;
		15'h3aa1: char_row_bitmap <= 16'b1111111111111100;
		15'h3aa2: char_row_bitmap <= 16'b1111111111111100;
		15'h3aa3: char_row_bitmap <= 16'b1111111111111100;
		15'h3aa4: char_row_bitmap <= 16'b1111111111111100;
		15'h3aa5: char_row_bitmap <= 16'b1111111111111100;
		15'h3aa6: char_row_bitmap <= 16'b1111111111111100;
		15'h3aa7: char_row_bitmap <= 16'b1111111111111100;
		15'h3aa8: char_row_bitmap <= 16'b1111111111111100;
		15'h3aa9: char_row_bitmap <= 16'b1111111111111100;
		15'h3aaa: char_row_bitmap <= 16'b0000000000000000;
		15'h3aab: char_row_bitmap <= 16'b0000000000000000;
		15'h3aac: char_row_bitmap <= 16'b1111111111111111;
		15'h3aad: char_row_bitmap <= 16'b1111111111111111;
		15'h3aae: char_row_bitmap <= 16'b1111111111111111;
		15'h3aaf: char_row_bitmap <= 16'b1111111111111111;
		15'h3ab0: char_row_bitmap <= 16'b1111111111111111;
		15'h3ab1: char_row_bitmap <= 16'b1111111111111111;
		15'h3ab2: char_row_bitmap <= 16'b1111111111111111;
		15'h3ab3: char_row_bitmap <= 16'b1111111111111111;
		15'h3ab4: char_row_bitmap <= 16'b1111111111111111;
		15'h3ab5: char_row_bitmap <= 16'b1111111111111111;
		15'h3ab6: char_row_bitmap <= 16'b1111111111111111;
		15'h3ab7: char_row_bitmap <= 16'b1111111111111111;
		15'h3ab8: char_row_bitmap <= 16'b1111111111111111;
		15'h3ab9: char_row_bitmap <= 16'b1111111111111111;
		15'h3aba: char_row_bitmap <= 16'b1111111111111111;
		15'h3abb: char_row_bitmap <= 16'b1111111111111111;
		15'h3abc: char_row_bitmap <= 16'b1111111111111111;
		15'h3abd: char_row_bitmap <= 16'b1111111111111111;
		15'h3abe: char_row_bitmap <= 16'b0000000000000000;
		15'h3abf: char_row_bitmap <= 16'b0000000000000000;
		15'h3ac0: char_row_bitmap <= 16'b0000000000000011;
		15'h3ac1: char_row_bitmap <= 16'b0000000000000011;
		15'h3ac2: char_row_bitmap <= 16'b0000000000000011;
		15'h3ac3: char_row_bitmap <= 16'b0000000000000011;
		15'h3ac4: char_row_bitmap <= 16'b0000000000000011;
		15'h3ac5: char_row_bitmap <= 16'b0000000000000011;
		15'h3ac6: char_row_bitmap <= 16'b0000000000000011;
		15'h3ac7: char_row_bitmap <= 16'b0000000000000011;
		15'h3ac8: char_row_bitmap <= 16'b0000000000000011;
		15'h3ac9: char_row_bitmap <= 16'b0000000000000011;
		15'h3aca: char_row_bitmap <= 16'b0000000000000011;
		15'h3acb: char_row_bitmap <= 16'b0000000000000011;
		15'h3acc: char_row_bitmap <= 16'b0000000000000011;
		15'h3acd: char_row_bitmap <= 16'b0000000000000011;
		15'h3ace: char_row_bitmap <= 16'b0000000000000011;
		15'h3acf: char_row_bitmap <= 16'b0000000000000011;
		15'h3ad0: char_row_bitmap <= 16'b0000000000000011;
		15'h3ad1: char_row_bitmap <= 16'b0000000000000011;
		15'h3ad2: char_row_bitmap <= 16'b0000000000000011;
		15'h3ad3: char_row_bitmap <= 16'b0000000000000011;
		15'h3ad4: char_row_bitmap <= 16'b0000000000001111;
		15'h3ad5: char_row_bitmap <= 16'b0000000000001111;
		15'h3ad6: char_row_bitmap <= 16'b0000000000001111;
		15'h3ad7: char_row_bitmap <= 16'b0000000000001111;
		15'h3ad8: char_row_bitmap <= 16'b0000000000001111;
		15'h3ad9: char_row_bitmap <= 16'b0000000000001111;
		15'h3ada: char_row_bitmap <= 16'b0000000000001111;
		15'h3adb: char_row_bitmap <= 16'b0000000000001111;
		15'h3adc: char_row_bitmap <= 16'b0000000000001111;
		15'h3add: char_row_bitmap <= 16'b0000000000001111;
		15'h3ade: char_row_bitmap <= 16'b0000000000001111;
		15'h3adf: char_row_bitmap <= 16'b0000000000001111;
		15'h3ae0: char_row_bitmap <= 16'b0000000000001111;
		15'h3ae1: char_row_bitmap <= 16'b0000000000001111;
		15'h3ae2: char_row_bitmap <= 16'b0000000000001111;
		15'h3ae3: char_row_bitmap <= 16'b0000000000001111;
		15'h3ae4: char_row_bitmap <= 16'b0000000000001111;
		15'h3ae5: char_row_bitmap <= 16'b0000000000001111;
		15'h3ae6: char_row_bitmap <= 16'b0000000000001111;
		15'h3ae7: char_row_bitmap <= 16'b0000000000001111;
		15'h3ae8: char_row_bitmap <= 16'b0000000000111111;
		15'h3ae9: char_row_bitmap <= 16'b0000000000111111;
		15'h3aea: char_row_bitmap <= 16'b0000000000111111;
		15'h3aeb: char_row_bitmap <= 16'b0000000000111111;
		15'h3aec: char_row_bitmap <= 16'b0000000000111111;
		15'h3aed: char_row_bitmap <= 16'b0000000000111111;
		15'h3aee: char_row_bitmap <= 16'b0000000000111111;
		15'h3aef: char_row_bitmap <= 16'b0000000000111111;
		15'h3af0: char_row_bitmap <= 16'b0000000000111111;
		15'h3af1: char_row_bitmap <= 16'b0000000000111111;
		15'h3af2: char_row_bitmap <= 16'b0000000000111111;
		15'h3af3: char_row_bitmap <= 16'b0000000000111111;
		15'h3af4: char_row_bitmap <= 16'b0000000000111111;
		15'h3af5: char_row_bitmap <= 16'b0000000000111111;
		15'h3af6: char_row_bitmap <= 16'b0000000000111111;
		15'h3af7: char_row_bitmap <= 16'b0000000000111111;
		15'h3af8: char_row_bitmap <= 16'b0000000000111111;
		15'h3af9: char_row_bitmap <= 16'b0000000000111111;
		15'h3afa: char_row_bitmap <= 16'b0000000000111111;
		15'h3afb: char_row_bitmap <= 16'b0000000000111111;
		15'h3afc: char_row_bitmap <= 16'b0000000011111111;
		15'h3afd: char_row_bitmap <= 16'b0000000011111111;
		15'h3afe: char_row_bitmap <= 16'b0000000011111111;
		15'h3aff: char_row_bitmap <= 16'b0000000011111111;
		15'h3b00: char_row_bitmap <= 16'b0000000011111111;
		15'h3b01: char_row_bitmap <= 16'b0000000011111111;
		15'h3b02: char_row_bitmap <= 16'b0000000011111111;
		15'h3b03: char_row_bitmap <= 16'b0000000011111111;
		15'h3b04: char_row_bitmap <= 16'b0000000011111111;
		15'h3b05: char_row_bitmap <= 16'b0000000011111111;
		15'h3b06: char_row_bitmap <= 16'b0000000011111111;
		15'h3b07: char_row_bitmap <= 16'b0000000011111111;
		15'h3b08: char_row_bitmap <= 16'b0000000011111111;
		15'h3b09: char_row_bitmap <= 16'b0000000011111111;
		15'h3b0a: char_row_bitmap <= 16'b0000000011111111;
		15'h3b0b: char_row_bitmap <= 16'b0000000011111111;
		15'h3b0c: char_row_bitmap <= 16'b0000000011111111;
		15'h3b0d: char_row_bitmap <= 16'b0000000011111111;
		15'h3b0e: char_row_bitmap <= 16'b0000000011111111;
		15'h3b0f: char_row_bitmap <= 16'b0000000011111111;
		15'h3b10: char_row_bitmap <= 16'b0000001111111111;
		15'h3b11: char_row_bitmap <= 16'b0000001111111111;
		15'h3b12: char_row_bitmap <= 16'b0000001111111111;
		15'h3b13: char_row_bitmap <= 16'b0000001111111111;
		15'h3b14: char_row_bitmap <= 16'b0000001111111111;
		15'h3b15: char_row_bitmap <= 16'b0000001111111111;
		15'h3b16: char_row_bitmap <= 16'b0000001111111111;
		15'h3b17: char_row_bitmap <= 16'b0000001111111111;
		15'h3b18: char_row_bitmap <= 16'b0000001111111111;
		15'h3b19: char_row_bitmap <= 16'b0000001111111111;
		15'h3b1a: char_row_bitmap <= 16'b0000001111111111;
		15'h3b1b: char_row_bitmap <= 16'b0000001111111111;
		15'h3b1c: char_row_bitmap <= 16'b0000001111111111;
		15'h3b1d: char_row_bitmap <= 16'b0000001111111111;
		15'h3b1e: char_row_bitmap <= 16'b0000001111111111;
		15'h3b1f: char_row_bitmap <= 16'b0000001111111111;
		15'h3b20: char_row_bitmap <= 16'b0000001111111111;
		15'h3b21: char_row_bitmap <= 16'b0000001111111111;
		15'h3b22: char_row_bitmap <= 16'b0000001111111111;
		15'h3b23: char_row_bitmap <= 16'b0000001111111111;
		15'h3b24: char_row_bitmap <= 16'b0000111111111111;
		15'h3b25: char_row_bitmap <= 16'b0000111111111111;
		15'h3b26: char_row_bitmap <= 16'b0000111111111111;
		15'h3b27: char_row_bitmap <= 16'b0000111111111111;
		15'h3b28: char_row_bitmap <= 16'b0000111111111111;
		15'h3b29: char_row_bitmap <= 16'b0000111111111111;
		15'h3b2a: char_row_bitmap <= 16'b0000111111111111;
		15'h3b2b: char_row_bitmap <= 16'b0000111111111111;
		15'h3b2c: char_row_bitmap <= 16'b0000111111111111;
		15'h3b2d: char_row_bitmap <= 16'b0000111111111111;
		15'h3b2e: char_row_bitmap <= 16'b0000111111111111;
		15'h3b2f: char_row_bitmap <= 16'b0000111111111111;
		15'h3b30: char_row_bitmap <= 16'b0000111111111111;
		15'h3b31: char_row_bitmap <= 16'b0000111111111111;
		15'h3b32: char_row_bitmap <= 16'b0000111111111111;
		15'h3b33: char_row_bitmap <= 16'b0000111111111111;
		15'h3b34: char_row_bitmap <= 16'b0000111111111111;
		15'h3b35: char_row_bitmap <= 16'b0000111111111111;
		15'h3b36: char_row_bitmap <= 16'b0000111111111111;
		15'h3b37: char_row_bitmap <= 16'b0000111111111111;
		15'h3b38: char_row_bitmap <= 16'b0011111111111111;
		15'h3b39: char_row_bitmap <= 16'b0011111111111111;
		15'h3b3a: char_row_bitmap <= 16'b0011111111111111;
		15'h3b3b: char_row_bitmap <= 16'b0011111111111111;
		15'h3b3c: char_row_bitmap <= 16'b0011111111111111;
		15'h3b3d: char_row_bitmap <= 16'b0011111111111111;
		15'h3b3e: char_row_bitmap <= 16'b0011111111111111;
		15'h3b3f: char_row_bitmap <= 16'b0011111111111111;
		15'h3b40: char_row_bitmap <= 16'b0011111111111111;
		15'h3b41: char_row_bitmap <= 16'b0011111111111111;
		15'h3b42: char_row_bitmap <= 16'b0011111111111111;
		15'h3b43: char_row_bitmap <= 16'b0011111111111111;
		15'h3b44: char_row_bitmap <= 16'b0011111111111111;
		15'h3b45: char_row_bitmap <= 16'b0011111111111111;
		15'h3b46: char_row_bitmap <= 16'b0011111111111111;
		15'h3b47: char_row_bitmap <= 16'b0011111111111111;
		15'h3b48: char_row_bitmap <= 16'b0011111111111111;
		15'h3b49: char_row_bitmap <= 16'b0011111111111111;
		15'h3b4a: char_row_bitmap <= 16'b0011111111111111;
		15'h3b4b: char_row_bitmap <= 16'b0011111111111111;
		15'h3b4c: char_row_bitmap <= 16'b1111111111111111;
		15'h3b4d: char_row_bitmap <= 16'b1111111111111111;
		15'h3b4e: char_row_bitmap <= 16'b1111111111111111;
		15'h3b4f: char_row_bitmap <= 16'b1111111111111111;
		15'h3b50: char_row_bitmap <= 16'b1111111111111111;
		15'h3b51: char_row_bitmap <= 16'b1111111111111111;
		15'h3b52: char_row_bitmap <= 16'b1111111111111111;
		15'h3b53: char_row_bitmap <= 16'b1111111111111111;
		15'h3b54: char_row_bitmap <= 16'b1111111111111111;
		15'h3b55: char_row_bitmap <= 16'b1111111111111111;
		15'h3b56: char_row_bitmap <= 16'b1111111111111111;
		15'h3b57: char_row_bitmap <= 16'b1111111111111111;
		15'h3b58: char_row_bitmap <= 16'b1111111111111111;
		15'h3b59: char_row_bitmap <= 16'b1111111111111111;
		15'h3b5a: char_row_bitmap <= 16'b1111111111111111;
		15'h3b5b: char_row_bitmap <= 16'b1111111111111111;
		15'h3b5c: char_row_bitmap <= 16'b1111111111111111;
		15'h3b5d: char_row_bitmap <= 16'b1111111111111111;
		15'h3b5e: char_row_bitmap <= 16'b1111111111111111;
		15'h3b5f: char_row_bitmap <= 16'b1111111111111111;
		15'h3b60: char_row_bitmap <= 16'b0000000000000001;
		15'h3b61: char_row_bitmap <= 16'b0000000000000001;
		15'h3b62: char_row_bitmap <= 16'b0000000000000001;
		15'h3b63: char_row_bitmap <= 16'b0000000000000001;
		15'h3b64: char_row_bitmap <= 16'b0000000000000001;
		15'h3b65: char_row_bitmap <= 16'b0000000000000001;
		15'h3b66: char_row_bitmap <= 16'b0000000000000001;
		15'h3b67: char_row_bitmap <= 16'b0000000000000001;
		15'h3b68: char_row_bitmap <= 16'b0000000000000001;
		15'h3b69: char_row_bitmap <= 16'b0000000000000001;
		15'h3b6a: char_row_bitmap <= 16'b0000000000000001;
		15'h3b6b: char_row_bitmap <= 16'b0000000000000001;
		15'h3b6c: char_row_bitmap <= 16'b0000000000000001;
		15'h3b6d: char_row_bitmap <= 16'b0000000000000001;
		15'h3b6e: char_row_bitmap <= 16'b0000000000000001;
		15'h3b6f: char_row_bitmap <= 16'b0000000000000001;
		15'h3b70: char_row_bitmap <= 16'b0000000000000001;
		15'h3b71: char_row_bitmap <= 16'b0000000000000001;
		15'h3b72: char_row_bitmap <= 16'b0000000000000000;
		15'h3b73: char_row_bitmap <= 16'b0000000000000000;
		15'h3b74: char_row_bitmap <= 16'b0000000000001111;
		15'h3b75: char_row_bitmap <= 16'b0000000000001111;
		15'h3b76: char_row_bitmap <= 16'b0000000000001111;
		15'h3b77: char_row_bitmap <= 16'b0000000000001111;
		15'h3b78: char_row_bitmap <= 16'b0000000000001111;
		15'h3b79: char_row_bitmap <= 16'b0000000000001111;
		15'h3b7a: char_row_bitmap <= 16'b0000000000001111;
		15'h3b7b: char_row_bitmap <= 16'b0000000000001111;
		15'h3b7c: char_row_bitmap <= 16'b0000000000001111;
		15'h3b7d: char_row_bitmap <= 16'b0000000000001111;
		15'h3b7e: char_row_bitmap <= 16'b0000000000001111;
		15'h3b7f: char_row_bitmap <= 16'b0000000000001111;
		15'h3b80: char_row_bitmap <= 16'b0000000000001111;
		15'h3b81: char_row_bitmap <= 16'b0000000000001111;
		15'h3b82: char_row_bitmap <= 16'b0000000000001111;
		15'h3b83: char_row_bitmap <= 16'b0000000000001111;
		15'h3b84: char_row_bitmap <= 16'b0000000000001111;
		15'h3b85: char_row_bitmap <= 16'b0000000000001111;
		15'h3b86: char_row_bitmap <= 16'b0000000000000000;
		15'h3b87: char_row_bitmap <= 16'b0000000000000000;
		15'h3b88: char_row_bitmap <= 16'b0000000000111111;
		15'h3b89: char_row_bitmap <= 16'b0000000000111111;
		15'h3b8a: char_row_bitmap <= 16'b0000000000111111;
		15'h3b8b: char_row_bitmap <= 16'b0000000000111111;
		15'h3b8c: char_row_bitmap <= 16'b0000000000111111;
		15'h3b8d: char_row_bitmap <= 16'b0000000000111111;
		15'h3b8e: char_row_bitmap <= 16'b0000000000111111;
		15'h3b8f: char_row_bitmap <= 16'b0000000000111111;
		15'h3b90: char_row_bitmap <= 16'b0000000000111111;
		15'h3b91: char_row_bitmap <= 16'b0000000000111111;
		15'h3b92: char_row_bitmap <= 16'b0000000000111111;
		15'h3b93: char_row_bitmap <= 16'b0000000000111111;
		15'h3b94: char_row_bitmap <= 16'b0000000000111111;
		15'h3b95: char_row_bitmap <= 16'b0000000000111111;
		15'h3b96: char_row_bitmap <= 16'b0000000000111111;
		15'h3b97: char_row_bitmap <= 16'b0000000000111111;
		15'h3b98: char_row_bitmap <= 16'b0000000000111111;
		15'h3b99: char_row_bitmap <= 16'b0000000000111111;
		15'h3b9a: char_row_bitmap <= 16'b0000000000000000;
		15'h3b9b: char_row_bitmap <= 16'b0000000000000000;
		15'h3b9c: char_row_bitmap <= 16'b0000000011111111;
		15'h3b9d: char_row_bitmap <= 16'b0000000011111111;
		15'h3b9e: char_row_bitmap <= 16'b0000000011111111;
		15'h3b9f: char_row_bitmap <= 16'b0000000011111111;
		15'h3ba0: char_row_bitmap <= 16'b0000000011111111;
		15'h3ba1: char_row_bitmap <= 16'b0000000011111111;
		15'h3ba2: char_row_bitmap <= 16'b0000000011111111;
		15'h3ba3: char_row_bitmap <= 16'b0000000011111111;
		15'h3ba4: char_row_bitmap <= 16'b0000000011111111;
		15'h3ba5: char_row_bitmap <= 16'b0000000011111111;
		15'h3ba6: char_row_bitmap <= 16'b0000000011111111;
		15'h3ba7: char_row_bitmap <= 16'b0000000011111111;
		15'h3ba8: char_row_bitmap <= 16'b0000000011111111;
		15'h3ba9: char_row_bitmap <= 16'b0000000011111111;
		15'h3baa: char_row_bitmap <= 16'b0000000011111111;
		15'h3bab: char_row_bitmap <= 16'b0000000011111111;
		15'h3bac: char_row_bitmap <= 16'b0000000011111111;
		15'h3bad: char_row_bitmap <= 16'b0000000011111111;
		15'h3bae: char_row_bitmap <= 16'b0000000000000000;
		15'h3baf: char_row_bitmap <= 16'b0000000000000000;
		15'h3bb0: char_row_bitmap <= 16'b0000001111111111;
		15'h3bb1: char_row_bitmap <= 16'b0000001111111111;
		15'h3bb2: char_row_bitmap <= 16'b0000001111111111;
		15'h3bb3: char_row_bitmap <= 16'b0000001111111111;
		15'h3bb4: char_row_bitmap <= 16'b0000001111111111;
		15'h3bb5: char_row_bitmap <= 16'b0000001111111111;
		15'h3bb6: char_row_bitmap <= 16'b0000001111111111;
		15'h3bb7: char_row_bitmap <= 16'b0000001111111111;
		15'h3bb8: char_row_bitmap <= 16'b0000001111111111;
		15'h3bb9: char_row_bitmap <= 16'b0000001111111111;
		15'h3bba: char_row_bitmap <= 16'b0000001111111111;
		15'h3bbb: char_row_bitmap <= 16'b0000001111111111;
		15'h3bbc: char_row_bitmap <= 16'b0000001111111111;
		15'h3bbd: char_row_bitmap <= 16'b0000001111111111;
		15'h3bbe: char_row_bitmap <= 16'b0000001111111111;
		15'h3bbf: char_row_bitmap <= 16'b0000001111111111;
		15'h3bc0: char_row_bitmap <= 16'b0000001111111111;
		15'h3bc1: char_row_bitmap <= 16'b0000001111111111;
		15'h3bc2: char_row_bitmap <= 16'b0000000000000000;
		15'h3bc3: char_row_bitmap <= 16'b0000000000000000;
		15'h3bc4: char_row_bitmap <= 16'b0000111111111111;
		15'h3bc5: char_row_bitmap <= 16'b0000111111111111;
		15'h3bc6: char_row_bitmap <= 16'b0000111111111111;
		15'h3bc7: char_row_bitmap <= 16'b0000111111111111;
		15'h3bc8: char_row_bitmap <= 16'b0000111111111111;
		15'h3bc9: char_row_bitmap <= 16'b0000111111111111;
		15'h3bca: char_row_bitmap <= 16'b0000111111111111;
		15'h3bcb: char_row_bitmap <= 16'b0000111111111111;
		15'h3bcc: char_row_bitmap <= 16'b0000111111111111;
		15'h3bcd: char_row_bitmap <= 16'b0000111111111111;
		15'h3bce: char_row_bitmap <= 16'b0000111111111111;
		15'h3bcf: char_row_bitmap <= 16'b0000111111111111;
		15'h3bd0: char_row_bitmap <= 16'b0000111111111111;
		15'h3bd1: char_row_bitmap <= 16'b0000111111111111;
		15'h3bd2: char_row_bitmap <= 16'b0000111111111111;
		15'h3bd3: char_row_bitmap <= 16'b0000111111111111;
		15'h3bd4: char_row_bitmap <= 16'b0000111111111111;
		15'h3bd5: char_row_bitmap <= 16'b0000111111111111;
		15'h3bd6: char_row_bitmap <= 16'b0000000000000000;
		15'h3bd7: char_row_bitmap <= 16'b0000000000000000;
		15'h3bd8: char_row_bitmap <= 16'b0011111111111111;
		15'h3bd9: char_row_bitmap <= 16'b0011111111111111;
		15'h3bda: char_row_bitmap <= 16'b0011111111111111;
		15'h3bdb: char_row_bitmap <= 16'b0011111111111111;
		15'h3bdc: char_row_bitmap <= 16'b0011111111111111;
		15'h3bdd: char_row_bitmap <= 16'b0011111111111111;
		15'h3bde: char_row_bitmap <= 16'b0011111111111111;
		15'h3bdf: char_row_bitmap <= 16'b0011111111111111;
		15'h3be0: char_row_bitmap <= 16'b0011111111111111;
		15'h3be1: char_row_bitmap <= 16'b0011111111111111;
		15'h3be2: char_row_bitmap <= 16'b0011111111111111;
		15'h3be3: char_row_bitmap <= 16'b0011111111111111;
		15'h3be4: char_row_bitmap <= 16'b0011111111111111;
		15'h3be5: char_row_bitmap <= 16'b0011111111111111;
		15'h3be6: char_row_bitmap <= 16'b0011111111111111;
		15'h3be7: char_row_bitmap <= 16'b0011111111111111;
		15'h3be8: char_row_bitmap <= 16'b0011111111111111;
		15'h3be9: char_row_bitmap <= 16'b0011111111111111;
		15'h3bea: char_row_bitmap <= 16'b0000000000000000;
		15'h3beb: char_row_bitmap <= 16'b0000000000000000;
		15'h3bec: char_row_bitmap <= 16'b1111111111111111;
		15'h3bed: char_row_bitmap <= 16'b1111111111111111;
		15'h3bee: char_row_bitmap <= 16'b1111111111111111;
		15'h3bef: char_row_bitmap <= 16'b1111111111111111;
		15'h3bf0: char_row_bitmap <= 16'b1111111111111111;
		15'h3bf1: char_row_bitmap <= 16'b1111111111111111;
		15'h3bf2: char_row_bitmap <= 16'b1111111111111111;
		15'h3bf3: char_row_bitmap <= 16'b1111111111111111;
		15'h3bf4: char_row_bitmap <= 16'b1111111111111111;
		15'h3bf5: char_row_bitmap <= 16'b1111111111111111;
		15'h3bf6: char_row_bitmap <= 16'b1111111111111111;
		15'h3bf7: char_row_bitmap <= 16'b1111111111111111;
		15'h3bf8: char_row_bitmap <= 16'b1111111111111111;
		15'h3bf9: char_row_bitmap <= 16'b1111111111111111;
		15'h3bfa: char_row_bitmap <= 16'b1111111111111111;
		15'h3bfb: char_row_bitmap <= 16'b1111111111111111;
		15'h3bfc: char_row_bitmap <= 16'b1111111111111111;
		15'h3bfd: char_row_bitmap <= 16'b1111111111111111;
		15'h3bfe: char_row_bitmap <= 16'b0000000000000000;
		15'h3bff: char_row_bitmap <= 16'b0000000000000000;
		15'h3c00: char_row_bitmap <= 16'b0000000000000000;
		15'h3c01: char_row_bitmap <= 16'b0000000000000000;
		15'h3c02: char_row_bitmap <= 16'b0000000000000000;
		15'h3c03: char_row_bitmap <= 16'b0000000000000000;
		15'h3c04: char_row_bitmap <= 16'b0000000000000000;
		15'h3c05: char_row_bitmap <= 16'b0000000000000000;
		15'h3c06: char_row_bitmap <= 16'b0000000000000000;
		15'h3c07: char_row_bitmap <= 16'b0000000000000000;
		15'h3c08: char_row_bitmap <= 16'b0000000000000000;
		15'h3c09: char_row_bitmap <= 16'b0000000000000000;
		15'h3c0a: char_row_bitmap <= 16'b0000000000000000;
		15'h3c0b: char_row_bitmap <= 16'b0000000000000000;
		15'h3c0c: char_row_bitmap <= 16'b0000000000000000;
		15'h3c0d: char_row_bitmap <= 16'b0000000000000000;
		15'h3c0e: char_row_bitmap <= 16'b0000000000000000;
		15'h3c0f: char_row_bitmap <= 16'b0000000000000000;
		15'h3c10: char_row_bitmap <= 16'b0000000000000000;
		15'h3c11: char_row_bitmap <= 16'b0000000000000000;
		15'h3c12: char_row_bitmap <= 16'b1111111111111111;
		15'h3c13: char_row_bitmap <= 16'b1111111111111111;
		15'h3c14: char_row_bitmap <= 16'b0000000000000000;
		15'h3c15: char_row_bitmap <= 16'b0000000000000000;
		15'h3c16: char_row_bitmap <= 16'b0000000000000000;
		15'h3c17: char_row_bitmap <= 16'b0000000000000000;
		15'h3c18: char_row_bitmap <= 16'b0000000000000000;
		15'h3c19: char_row_bitmap <= 16'b0000000000000000;
		15'h3c1a: char_row_bitmap <= 16'b0000000000000000;
		15'h3c1b: char_row_bitmap <= 16'b0000000000000000;
		15'h3c1c: char_row_bitmap <= 16'b0000000000000000;
		15'h3c1d: char_row_bitmap <= 16'b0000000000000000;
		15'h3c1e: char_row_bitmap <= 16'b0000000000000000;
		15'h3c1f: char_row_bitmap <= 16'b0000000000000000;
		15'h3c20: char_row_bitmap <= 16'b0000000000000000;
		15'h3c21: char_row_bitmap <= 16'b0000000000000000;
		15'h3c22: char_row_bitmap <= 16'b0000000000000000;
		15'h3c23: char_row_bitmap <= 16'b0000000000000000;
		15'h3c24: char_row_bitmap <= 16'b1111111111111111;
		15'h3c25: char_row_bitmap <= 16'b1111111111111111;
		15'h3c26: char_row_bitmap <= 16'b1111111111111111;
		15'h3c27: char_row_bitmap <= 16'b1111111111111111;
		15'h3c28: char_row_bitmap <= 16'b0000000000000000;
		15'h3c29: char_row_bitmap <= 16'b0000000000000000;
		15'h3c2a: char_row_bitmap <= 16'b0000000000000000;
		15'h3c2b: char_row_bitmap <= 16'b0000000000000000;
		15'h3c2c: char_row_bitmap <= 16'b0000000000000000;
		15'h3c2d: char_row_bitmap <= 16'b0000000000000000;
		15'h3c2e: char_row_bitmap <= 16'b0000000000000000;
		15'h3c2f: char_row_bitmap <= 16'b0000000000000000;
		15'h3c30: char_row_bitmap <= 16'b0000000000000000;
		15'h3c31: char_row_bitmap <= 16'b0000000000000000;
		15'h3c32: char_row_bitmap <= 16'b0000000000000000;
		15'h3c33: char_row_bitmap <= 16'b0000000000000000;
		15'h3c34: char_row_bitmap <= 16'b0000000000000000;
		15'h3c35: char_row_bitmap <= 16'b0000000000000000;
		15'h3c36: char_row_bitmap <= 16'b1111111111111111;
		15'h3c37: char_row_bitmap <= 16'b1111111111111111;
		15'h3c38: char_row_bitmap <= 16'b1111111111111111;
		15'h3c39: char_row_bitmap <= 16'b1111111111111111;
		15'h3c3a: char_row_bitmap <= 16'b1111111111111111;
		15'h3c3b: char_row_bitmap <= 16'b1111111111111111;
		15'h3c3c: char_row_bitmap <= 16'b0000000000000000;
		15'h3c3d: char_row_bitmap <= 16'b0000000000000000;
		15'h3c3e: char_row_bitmap <= 16'b0000000000000000;
		15'h3c3f: char_row_bitmap <= 16'b0000000000000000;
		15'h3c40: char_row_bitmap <= 16'b0000000000000000;
		15'h3c41: char_row_bitmap <= 16'b0000000000000000;
		15'h3c42: char_row_bitmap <= 16'b0000000000000000;
		15'h3c43: char_row_bitmap <= 16'b0000000000000000;
		15'h3c44: char_row_bitmap <= 16'b0000000000000000;
		15'h3c45: char_row_bitmap <= 16'b0000000000000000;
		15'h3c46: char_row_bitmap <= 16'b0000000000000000;
		15'h3c47: char_row_bitmap <= 16'b0000000000000000;
		15'h3c48: char_row_bitmap <= 16'b1111111111111111;
		15'h3c49: char_row_bitmap <= 16'b1111111111111111;
		15'h3c4a: char_row_bitmap <= 16'b1111111111111111;
		15'h3c4b: char_row_bitmap <= 16'b1111111111111111;
		15'h3c4c: char_row_bitmap <= 16'b1111111111111111;
		15'h3c4d: char_row_bitmap <= 16'b1111111111111111;
		15'h3c4e: char_row_bitmap <= 16'b1111111111111111;
		15'h3c4f: char_row_bitmap <= 16'b1111111111111111;
		15'h3c50: char_row_bitmap <= 16'b0000000000000000;
		15'h3c51: char_row_bitmap <= 16'b0000000000000000;
		15'h3c52: char_row_bitmap <= 16'b0000000000000000;
		15'h3c53: char_row_bitmap <= 16'b0000000000000000;
		15'h3c54: char_row_bitmap <= 16'b0000000000000000;
		15'h3c55: char_row_bitmap <= 16'b0000000000000000;
		15'h3c56: char_row_bitmap <= 16'b0000000000000000;
		15'h3c57: char_row_bitmap <= 16'b0000000000000000;
		15'h3c58: char_row_bitmap <= 16'b0000000000000000;
		15'h3c59: char_row_bitmap <= 16'b0000000000000000;
		15'h3c5a: char_row_bitmap <= 16'b1111111111111111;
		15'h3c5b: char_row_bitmap <= 16'b1111111111111111;
		15'h3c5c: char_row_bitmap <= 16'b1111111111111111;
		15'h3c5d: char_row_bitmap <= 16'b1111111111111111;
		15'h3c5e: char_row_bitmap <= 16'b1111111111111111;
		15'h3c5f: char_row_bitmap <= 16'b1111111111111111;
		15'h3c60: char_row_bitmap <= 16'b1111111111111111;
		15'h3c61: char_row_bitmap <= 16'b1111111111111111;
		15'h3c62: char_row_bitmap <= 16'b1111111111111111;
		15'h3c63: char_row_bitmap <= 16'b1111111111111111;
		15'h3c64: char_row_bitmap <= 16'b0000000000000000;
		15'h3c65: char_row_bitmap <= 16'b0000000000000000;
		15'h3c66: char_row_bitmap <= 16'b0000000000000000;
		15'h3c67: char_row_bitmap <= 16'b0000000000000000;
		15'h3c68: char_row_bitmap <= 16'b0000000000000000;
		15'h3c69: char_row_bitmap <= 16'b0000000000000000;
		15'h3c6a: char_row_bitmap <= 16'b0000000000000000;
		15'h3c6b: char_row_bitmap <= 16'b0000000000000000;
		15'h3c6c: char_row_bitmap <= 16'b1111111111111111;
		15'h3c6d: char_row_bitmap <= 16'b1111111111111111;
		15'h3c6e: char_row_bitmap <= 16'b1111111111111111;
		15'h3c6f: char_row_bitmap <= 16'b1111111111111111;
		15'h3c70: char_row_bitmap <= 16'b1111111111111111;
		15'h3c71: char_row_bitmap <= 16'b1111111111111111;
		15'h3c72: char_row_bitmap <= 16'b1111111111111111;
		15'h3c73: char_row_bitmap <= 16'b1111111111111111;
		15'h3c74: char_row_bitmap <= 16'b1111111111111111;
		15'h3c75: char_row_bitmap <= 16'b1111111111111111;
		15'h3c76: char_row_bitmap <= 16'b1111111111111111;
		15'h3c77: char_row_bitmap <= 16'b1111111111111111;
		15'h3c78: char_row_bitmap <= 16'b0000000000000000;
		15'h3c79: char_row_bitmap <= 16'b0000000000000000;
		15'h3c7a: char_row_bitmap <= 16'b0000000000000000;
		15'h3c7b: char_row_bitmap <= 16'b0000000000000000;
		15'h3c7c: char_row_bitmap <= 16'b0000000000000000;
		15'h3c7d: char_row_bitmap <= 16'b0000000000000000;
		15'h3c7e: char_row_bitmap <= 16'b1111111111111111;
		15'h3c7f: char_row_bitmap <= 16'b1111111111111111;
		15'h3c80: char_row_bitmap <= 16'b1111111111111111;
		15'h3c81: char_row_bitmap <= 16'b1111111111111111;
		15'h3c82: char_row_bitmap <= 16'b1111111111111111;
		15'h3c83: char_row_bitmap <= 16'b1111111111111111;
		15'h3c84: char_row_bitmap <= 16'b1111111111111111;
		15'h3c85: char_row_bitmap <= 16'b1111111111111111;
		15'h3c86: char_row_bitmap <= 16'b1111111111111111;
		15'h3c87: char_row_bitmap <= 16'b1111111111111111;
		15'h3c88: char_row_bitmap <= 16'b1111111111111111;
		15'h3c89: char_row_bitmap <= 16'b1111111111111111;
		15'h3c8a: char_row_bitmap <= 16'b1111111111111111;
		15'h3c8b: char_row_bitmap <= 16'b1111111111111111;
		15'h3c8c: char_row_bitmap <= 16'b0000000000000000;
		15'h3c8d: char_row_bitmap <= 16'b0000000000000000;
		15'h3c8e: char_row_bitmap <= 16'b0000000000000000;
		15'h3c8f: char_row_bitmap <= 16'b0000000000000000;
		15'h3c90: char_row_bitmap <= 16'b1111111111111111;
		15'h3c91: char_row_bitmap <= 16'b1111111111111111;
		15'h3c92: char_row_bitmap <= 16'b1111111111111111;
		15'h3c93: char_row_bitmap <= 16'b1111111111111111;
		15'h3c94: char_row_bitmap <= 16'b1111111111111111;
		15'h3c95: char_row_bitmap <= 16'b1111111111111111;
		15'h3c96: char_row_bitmap <= 16'b1111111111111111;
		15'h3c97: char_row_bitmap <= 16'b1111111111111111;
		15'h3c98: char_row_bitmap <= 16'b1111111111111111;
		15'h3c99: char_row_bitmap <= 16'b1111111111111111;
		15'h3c9a: char_row_bitmap <= 16'b1111111111111111;
		15'h3c9b: char_row_bitmap <= 16'b1111111111111111;
		15'h3c9c: char_row_bitmap <= 16'b1111111111111111;
		15'h3c9d: char_row_bitmap <= 16'b1111111111111111;
		15'h3c9e: char_row_bitmap <= 16'b1111111111111111;
		15'h3c9f: char_row_bitmap <= 16'b1111111111111111;
		15'h3ca0: char_row_bitmap <= 16'b0000000000000000;
		15'h3ca1: char_row_bitmap <= 16'b0000000000000000;
		15'h3ca2: char_row_bitmap <= 16'b1111111111111111;
		15'h3ca3: char_row_bitmap <= 16'b1111111111111111;
		15'h3ca4: char_row_bitmap <= 16'b1111111111111111;
		15'h3ca5: char_row_bitmap <= 16'b1111111111111111;
		15'h3ca6: char_row_bitmap <= 16'b1111111111111111;
		15'h3ca7: char_row_bitmap <= 16'b1111111111111111;
		15'h3ca8: char_row_bitmap <= 16'b1111111111111111;
		15'h3ca9: char_row_bitmap <= 16'b1111111111111111;
		15'h3caa: char_row_bitmap <= 16'b1111111111111111;
		15'h3cab: char_row_bitmap <= 16'b1111111111111111;
		15'h3cac: char_row_bitmap <= 16'b1111111111111111;
		15'h3cad: char_row_bitmap <= 16'b1111111111111111;
		15'h3cae: char_row_bitmap <= 16'b1111111111111111;
		15'h3caf: char_row_bitmap <= 16'b1111111111111111;
		15'h3cb0: char_row_bitmap <= 16'b1111111111111111;
		15'h3cb1: char_row_bitmap <= 16'b1111111111111111;
		15'h3cb2: char_row_bitmap <= 16'b1111111111111111;
		15'h3cb3: char_row_bitmap <= 16'b1111111111111111;
		15'h3cb4: char_row_bitmap <= 16'b1111111111111111;
		15'h3cb5: char_row_bitmap <= 16'b1111111111111111;
		15'h3cb6: char_row_bitmap <= 16'b1111111111111111;
		15'h3cb7: char_row_bitmap <= 16'b1111111111111111;
		15'h3cb8: char_row_bitmap <= 16'b1111111111111111;
		15'h3cb9: char_row_bitmap <= 16'b1111111111111111;
		15'h3cba: char_row_bitmap <= 16'b1111111111111111;
		15'h3cbb: char_row_bitmap <= 16'b1111111111111111;
		15'h3cbc: char_row_bitmap <= 16'b1111111111111111;
		15'h3cbd: char_row_bitmap <= 16'b1111111111111111;
		15'h3cbe: char_row_bitmap <= 16'b1111111111111111;
		15'h3cbf: char_row_bitmap <= 16'b1111111111111111;
		15'h3cc0: char_row_bitmap <= 16'b1111111111111111;
		15'h3cc1: char_row_bitmap <= 16'b1111111111111111;
		15'h3cc2: char_row_bitmap <= 16'b1111111111111111;
		15'h3cc3: char_row_bitmap <= 16'b1111111111111111;
		15'h3cc4: char_row_bitmap <= 16'b1111111111111111;
		15'h3cc5: char_row_bitmap <= 16'b1111111111111111;
		15'h3cc6: char_row_bitmap <= 16'b1111111111111111;
		15'h3cc7: char_row_bitmap <= 16'b1111111111111111;
		15'h3cc8: char_row_bitmap <= 16'b1111111111111111;
		15'h3cc9: char_row_bitmap <= 16'b1111111111111111;
		15'h3cca: char_row_bitmap <= 16'b0000000000000011;
		15'h3ccb: char_row_bitmap <= 16'b0000000000000011;
		15'h3ccc: char_row_bitmap <= 16'b0000000000000011;
		15'h3ccd: char_row_bitmap <= 16'b0000000000000011;
		15'h3cce: char_row_bitmap <= 16'b0000000000000011;
		15'h3ccf: char_row_bitmap <= 16'b0000000000000011;
		15'h3cd0: char_row_bitmap <= 16'b0000000000000011;
		15'h3cd1: char_row_bitmap <= 16'b0000000000000011;
		15'h3cd2: char_row_bitmap <= 16'b0000000000000011;
		15'h3cd3: char_row_bitmap <= 16'b0000000000000011;
		15'h3cd4: char_row_bitmap <= 16'b0000000000000011;
		15'h3cd5: char_row_bitmap <= 16'b0000000000000011;
		15'h3cd6: char_row_bitmap <= 16'b0000000000000011;
		15'h3cd7: char_row_bitmap <= 16'b0000000000000011;
		15'h3cd8: char_row_bitmap <= 16'b0000000000000011;
		15'h3cd9: char_row_bitmap <= 16'b0000000000000011;
		15'h3cda: char_row_bitmap <= 16'b0000000000000011;
		15'h3cdb: char_row_bitmap <= 16'b0000000000000011;
		15'h3cdc: char_row_bitmap <= 16'b0000000000000011;
		15'h3cdd: char_row_bitmap <= 16'b0000000000000011;
		15'h3cde: char_row_bitmap <= 16'b0000000000000011;
		15'h3cdf: char_row_bitmap <= 16'b0000000000000011;
		15'h3ce0: char_row_bitmap <= 16'b0000000000000011;
		15'h3ce1: char_row_bitmap <= 16'b0000000000000011;
		15'h3ce2: char_row_bitmap <= 16'b0000000000000011;
		15'h3ce3: char_row_bitmap <= 16'b0000000000000011;
		15'h3ce4: char_row_bitmap <= 16'b0000000000000011;
		15'h3ce5: char_row_bitmap <= 16'b0000000000000011;
		15'h3ce6: char_row_bitmap <= 16'b0000000000000011;
		15'h3ce7: char_row_bitmap <= 16'b0000000000000011;
		15'h3ce8: char_row_bitmap <= 16'b0000000000000011;
		15'h3ce9: char_row_bitmap <= 16'b0000000000000011;
		15'h3cea: char_row_bitmap <= 16'b0000000000000011;
		15'h3ceb: char_row_bitmap <= 16'b0000000000000011;
		15'h3cec: char_row_bitmap <= 16'b0000000000000011;
		15'h3ced: char_row_bitmap <= 16'b0000000000000011;
		15'h3cee: char_row_bitmap <= 16'b1111111111111111;
		15'h3cef: char_row_bitmap <= 16'b1111111111111111;
		15'h3cf0: char_row_bitmap <= 16'b1100000000000000;
		15'h3cf1: char_row_bitmap <= 16'b1100000000000000;
		15'h3cf2: char_row_bitmap <= 16'b1100000000000000;
		15'h3cf3: char_row_bitmap <= 16'b1100000000000000;
		15'h3cf4: char_row_bitmap <= 16'b1100000000000000;
		15'h3cf5: char_row_bitmap <= 16'b1100000000000000;
		15'h3cf6: char_row_bitmap <= 16'b1100000000000000;
		15'h3cf7: char_row_bitmap <= 16'b1100000000000000;
		15'h3cf8: char_row_bitmap <= 16'b1100000000000000;
		15'h3cf9: char_row_bitmap <= 16'b1100000000000000;
		15'h3cfa: char_row_bitmap <= 16'b1100000000000000;
		15'h3cfb: char_row_bitmap <= 16'b1100000000000000;
		15'h3cfc: char_row_bitmap <= 16'b1100000000000000;
		15'h3cfd: char_row_bitmap <= 16'b1100000000000000;
		15'h3cfe: char_row_bitmap <= 16'b1100000000000000;
		15'h3cff: char_row_bitmap <= 16'b1100000000000000;
		15'h3d00: char_row_bitmap <= 16'b1100000000000000;
		15'h3d01: char_row_bitmap <= 16'b1100000000000000;
		15'h3d02: char_row_bitmap <= 16'b1111111111111111;
		15'h3d03: char_row_bitmap <= 16'b1111111111111111;
		15'h3d04: char_row_bitmap <= 16'b1111111111111111;
		15'h3d05: char_row_bitmap <= 16'b1111111111111111;
		15'h3d06: char_row_bitmap <= 16'b1100000000000000;
		15'h3d07: char_row_bitmap <= 16'b1100000000000000;
		15'h3d08: char_row_bitmap <= 16'b1100000000000000;
		15'h3d09: char_row_bitmap <= 16'b1100000000000000;
		15'h3d0a: char_row_bitmap <= 16'b1100000000000000;
		15'h3d0b: char_row_bitmap <= 16'b1100000000000000;
		15'h3d0c: char_row_bitmap <= 16'b1100000000000000;
		15'h3d0d: char_row_bitmap <= 16'b1100000000000000;
		15'h3d0e: char_row_bitmap <= 16'b1100000000000000;
		15'h3d0f: char_row_bitmap <= 16'b1100000000000000;
		15'h3d10: char_row_bitmap <= 16'b1100000000000000;
		15'h3d11: char_row_bitmap <= 16'b1100000000000000;
		15'h3d12: char_row_bitmap <= 16'b1100000000000000;
		15'h3d13: char_row_bitmap <= 16'b1100000000000000;
		15'h3d14: char_row_bitmap <= 16'b1100000000000000;
		15'h3d15: char_row_bitmap <= 16'b1100000000000000;
		15'h3d16: char_row_bitmap <= 16'b1100000000000000;
		15'h3d17: char_row_bitmap <= 16'b1100000000000000;
		15'h3d18: char_row_bitmap <= 16'b1111111111111111;
		15'h3d19: char_row_bitmap <= 16'b1111111111111111;
		15'h3d1a: char_row_bitmap <= 16'b0000000000000000;
		15'h3d1b: char_row_bitmap <= 16'b0000000000000000;
		15'h3d1c: char_row_bitmap <= 16'b0000000000000000;
		15'h3d1d: char_row_bitmap <= 16'b0000000000000000;
		15'h3d1e: char_row_bitmap <= 16'b0000000000000000;
		15'h3d1f: char_row_bitmap <= 16'b0000000000000000;
		15'h3d20: char_row_bitmap <= 16'b0000000000000000;
		15'h3d21: char_row_bitmap <= 16'b0000000000000000;
		15'h3d22: char_row_bitmap <= 16'b0000000000000000;
		15'h3d23: char_row_bitmap <= 16'b0000000000000000;
		15'h3d24: char_row_bitmap <= 16'b0000000000000000;
		15'h3d25: char_row_bitmap <= 16'b0000000000000000;
		15'h3d26: char_row_bitmap <= 16'b0000000000000000;
		15'h3d27: char_row_bitmap <= 16'b0000000000000000;
		15'h3d28: char_row_bitmap <= 16'b0000000000000000;
		15'h3d29: char_row_bitmap <= 16'b0000000000000000;
		15'h3d2a: char_row_bitmap <= 16'b1111111111111111;
		15'h3d2b: char_row_bitmap <= 16'b1111111111111111;
		15'h3d2c: char_row_bitmap <= 16'b1100000000000011;
		15'h3d2d: char_row_bitmap <= 16'b1100000000000011;
		15'h3d2e: char_row_bitmap <= 16'b1100000000000011;
		15'h3d2f: char_row_bitmap <= 16'b1100000000000011;
		15'h3d30: char_row_bitmap <= 16'b1100000000000011;
		15'h3d31: char_row_bitmap <= 16'b1100000000000011;
		15'h3d32: char_row_bitmap <= 16'b1100000000000011;
		15'h3d33: char_row_bitmap <= 16'b1100000000000011;
		15'h3d34: char_row_bitmap <= 16'b1100000000000011;
		15'h3d35: char_row_bitmap <= 16'b1100000000000011;
		15'h3d36: char_row_bitmap <= 16'b1100000000000011;
		15'h3d37: char_row_bitmap <= 16'b1100000000000011;
		15'h3d38: char_row_bitmap <= 16'b1100000000000011;
		15'h3d39: char_row_bitmap <= 16'b1100000000000011;
		15'h3d3a: char_row_bitmap <= 16'b1100000000000011;
		15'h3d3b: char_row_bitmap <= 16'b1100000000000011;
		15'h3d3c: char_row_bitmap <= 16'b1100000000000011;
		15'h3d3d: char_row_bitmap <= 16'b1100000000000011;
		15'h3d3e: char_row_bitmap <= 16'b1100000000000011;
		15'h3d3f: char_row_bitmap <= 16'b1100000000000011;
		15'h3d40: char_row_bitmap <= 16'b0000000000000000;
		15'h3d41: char_row_bitmap <= 16'b0000000000000000;
		15'h3d42: char_row_bitmap <= 16'b0000000000000000;
		15'h3d43: char_row_bitmap <= 16'b0000000000000000;
		15'h3d44: char_row_bitmap <= 16'b0000000000000000;
		15'h3d45: char_row_bitmap <= 16'b0000000000000000;
		15'h3d46: char_row_bitmap <= 16'b0000000000000000;
		15'h3d47: char_row_bitmap <= 16'b0000000000000000;
		15'h3d48: char_row_bitmap <= 16'b0000000000000000;
		15'h3d49: char_row_bitmap <= 16'b0000000000000000;
		15'h3d4a: char_row_bitmap <= 16'b0000000000000000;
		15'h3d4b: char_row_bitmap <= 16'b0000000000000000;
		15'h3d4c: char_row_bitmap <= 16'b0000000000000000;
		15'h3d4d: char_row_bitmap <= 16'b0000000000000000;
		15'h3d4e: char_row_bitmap <= 16'b0000000000000000;
		15'h3d4f: char_row_bitmap <= 16'b0000000000000000;
		15'h3d50: char_row_bitmap <= 16'b0000000000000000;
		15'h3d51: char_row_bitmap <= 16'b0000000000000000;
		15'h3d52: char_row_bitmap <= 16'b1111111111111100;
		15'h3d53: char_row_bitmap <= 16'b1111111111111100;
		15'h3d54: char_row_bitmap <= 16'b0000000000000000;
		15'h3d55: char_row_bitmap <= 16'b0000000000000000;
		15'h3d56: char_row_bitmap <= 16'b0000000000000000;
		15'h3d57: char_row_bitmap <= 16'b0000000000000000;
		15'h3d58: char_row_bitmap <= 16'b0000000000000000;
		15'h3d59: char_row_bitmap <= 16'b0000000000000000;
		15'h3d5a: char_row_bitmap <= 16'b0000000000000000;
		15'h3d5b: char_row_bitmap <= 16'b0000000000000000;
		15'h3d5c: char_row_bitmap <= 16'b0000000000000000;
		15'h3d5d: char_row_bitmap <= 16'b0000000000000000;
		15'h3d5e: char_row_bitmap <= 16'b0000000000000000;
		15'h3d5f: char_row_bitmap <= 16'b0000000000000000;
		15'h3d60: char_row_bitmap <= 16'b0000000000000000;
		15'h3d61: char_row_bitmap <= 16'b0000000000000000;
		15'h3d62: char_row_bitmap <= 16'b0000000000000000;
		15'h3d63: char_row_bitmap <= 16'b0000000000000000;
		15'h3d64: char_row_bitmap <= 16'b1111111111111100;
		15'h3d65: char_row_bitmap <= 16'b1111111111111100;
		15'h3d66: char_row_bitmap <= 16'b1111111111111100;
		15'h3d67: char_row_bitmap <= 16'b1111111111111100;
		15'h3d68: char_row_bitmap <= 16'b0000000000000000;
		15'h3d69: char_row_bitmap <= 16'b0000000000000000;
		15'h3d6a: char_row_bitmap <= 16'b0000000000000000;
		15'h3d6b: char_row_bitmap <= 16'b0000000000000000;
		15'h3d6c: char_row_bitmap <= 16'b0000000000000000;
		15'h3d6d: char_row_bitmap <= 16'b0000000000000000;
		15'h3d6e: char_row_bitmap <= 16'b0000000000000000;
		15'h3d6f: char_row_bitmap <= 16'b0000000000000000;
		15'h3d70: char_row_bitmap <= 16'b0000000000000000;
		15'h3d71: char_row_bitmap <= 16'b0000000000000000;
		15'h3d72: char_row_bitmap <= 16'b0000000000000000;
		15'h3d73: char_row_bitmap <= 16'b0000000000000000;
		15'h3d74: char_row_bitmap <= 16'b0000000000000000;
		15'h3d75: char_row_bitmap <= 16'b0000000000000000;
		15'h3d76: char_row_bitmap <= 16'b1111111111111100;
		15'h3d77: char_row_bitmap <= 16'b1111111111111100;
		15'h3d78: char_row_bitmap <= 16'b1111111111111100;
		15'h3d79: char_row_bitmap <= 16'b1111111111111100;
		15'h3d7a: char_row_bitmap <= 16'b1111111111111100;
		15'h3d7b: char_row_bitmap <= 16'b1111111111111100;
		15'h3d7c: char_row_bitmap <= 16'b0000000000000000;
		15'h3d7d: char_row_bitmap <= 16'b0000000000000000;
		15'h3d7e: char_row_bitmap <= 16'b0000000000000000;
		15'h3d7f: char_row_bitmap <= 16'b0000000000000000;
		15'h3d80: char_row_bitmap <= 16'b0000000000000000;
		15'h3d81: char_row_bitmap <= 16'b0000000000000000;
		15'h3d82: char_row_bitmap <= 16'b0000000000000000;
		15'h3d83: char_row_bitmap <= 16'b0000000000000000;
		15'h3d84: char_row_bitmap <= 16'b0000000000000000;
		15'h3d85: char_row_bitmap <= 16'b0000000000000000;
		15'h3d86: char_row_bitmap <= 16'b0000000000000000;
		15'h3d87: char_row_bitmap <= 16'b0000000000000000;
		15'h3d88: char_row_bitmap <= 16'b1111111111111100;
		15'h3d89: char_row_bitmap <= 16'b1111111111111100;
		15'h3d8a: char_row_bitmap <= 16'b1111111111111100;
		15'h3d8b: char_row_bitmap <= 16'b1111111111111100;
		15'h3d8c: char_row_bitmap <= 16'b1111111111111100;
		15'h3d8d: char_row_bitmap <= 16'b1111111111111100;
		15'h3d8e: char_row_bitmap <= 16'b1111111111111100;
		15'h3d8f: char_row_bitmap <= 16'b1111111111111100;
		15'h3d90: char_row_bitmap <= 16'b0000000000000000;
		15'h3d91: char_row_bitmap <= 16'b0000000000000000;
		15'h3d92: char_row_bitmap <= 16'b0000000000000000;
		15'h3d93: char_row_bitmap <= 16'b0000000000000000;
		15'h3d94: char_row_bitmap <= 16'b0000000000000000;
		15'h3d95: char_row_bitmap <= 16'b0000000000000000;
		15'h3d96: char_row_bitmap <= 16'b0000000000000000;
		15'h3d97: char_row_bitmap <= 16'b0000000000000000;
		15'h3d98: char_row_bitmap <= 16'b0000000000000000;
		15'h3d99: char_row_bitmap <= 16'b0000000000000000;
		15'h3d9a: char_row_bitmap <= 16'b1111111111111100;
		15'h3d9b: char_row_bitmap <= 16'b1111111111111100;
		15'h3d9c: char_row_bitmap <= 16'b1111111111111100;
		15'h3d9d: char_row_bitmap <= 16'b1111111111111100;
		15'h3d9e: char_row_bitmap <= 16'b1111111111111100;
		15'h3d9f: char_row_bitmap <= 16'b1111111111111100;
		15'h3da0: char_row_bitmap <= 16'b1111111111111100;
		15'h3da1: char_row_bitmap <= 16'b1111111111111100;
		15'h3da2: char_row_bitmap <= 16'b1111111111111100;
		15'h3da3: char_row_bitmap <= 16'b1111111111111100;
		15'h3da4: char_row_bitmap <= 16'b0000000000000000;
		15'h3da5: char_row_bitmap <= 16'b0000000000000000;
		15'h3da6: char_row_bitmap <= 16'b0000000000000000;
		15'h3da7: char_row_bitmap <= 16'b0000000000000000;
		15'h3da8: char_row_bitmap <= 16'b0000000000000000;
		15'h3da9: char_row_bitmap <= 16'b0000000000000000;
		15'h3daa: char_row_bitmap <= 16'b0000000000000000;
		15'h3dab: char_row_bitmap <= 16'b0000000000000000;
		15'h3dac: char_row_bitmap <= 16'b1111111111111100;
		15'h3dad: char_row_bitmap <= 16'b1111111111111100;
		15'h3dae: char_row_bitmap <= 16'b1111111111111100;
		15'h3daf: char_row_bitmap <= 16'b1111111111111100;
		15'h3db0: char_row_bitmap <= 16'b1111111111111100;
		15'h3db1: char_row_bitmap <= 16'b1111111111111100;
		15'h3db2: char_row_bitmap <= 16'b1111111111111100;
		15'h3db3: char_row_bitmap <= 16'b1111111111111100;
		15'h3db4: char_row_bitmap <= 16'b1111111111111100;
		15'h3db5: char_row_bitmap <= 16'b1111111111111100;
		15'h3db6: char_row_bitmap <= 16'b1111111111111100;
		15'h3db7: char_row_bitmap <= 16'b1111111111111100;
		15'h3db8: char_row_bitmap <= 16'b0000000000000000;
		15'h3db9: char_row_bitmap <= 16'b0000000000000000;
		15'h3dba: char_row_bitmap <= 16'b0000000000000000;
		15'h3dbb: char_row_bitmap <= 16'b0000000000000000;
		15'h3dbc: char_row_bitmap <= 16'b0000000000000000;
		15'h3dbd: char_row_bitmap <= 16'b0000000000000000;
		15'h3dbe: char_row_bitmap <= 16'b1111111111111100;
		15'h3dbf: char_row_bitmap <= 16'b1111111111111100;
		15'h3dc0: char_row_bitmap <= 16'b1111111111111100;
		15'h3dc1: char_row_bitmap <= 16'b1111111111111100;
		15'h3dc2: char_row_bitmap <= 16'b1111111111111100;
		15'h3dc3: char_row_bitmap <= 16'b1111111111111100;
		15'h3dc4: char_row_bitmap <= 16'b1111111111111100;
		15'h3dc5: char_row_bitmap <= 16'b1111111111111100;
		15'h3dc6: char_row_bitmap <= 16'b1111111111111100;
		15'h3dc7: char_row_bitmap <= 16'b1111111111111100;
		15'h3dc8: char_row_bitmap <= 16'b1111111111111100;
		15'h3dc9: char_row_bitmap <= 16'b1111111111111100;
		15'h3dca: char_row_bitmap <= 16'b1111111111111100;
		15'h3dcb: char_row_bitmap <= 16'b1111111111111100;
		15'h3dcc: char_row_bitmap <= 16'b0000000000000000;
		15'h3dcd: char_row_bitmap <= 16'b0000000000000000;
		15'h3dce: char_row_bitmap <= 16'b0000000000000000;
		15'h3dcf: char_row_bitmap <= 16'b0000000000000000;
		15'h3dd0: char_row_bitmap <= 16'b1111111111111100;
		15'h3dd1: char_row_bitmap <= 16'b1111111111111100;
		15'h3dd2: char_row_bitmap <= 16'b1111111111111100;
		15'h3dd3: char_row_bitmap <= 16'b1111111111111100;
		15'h3dd4: char_row_bitmap <= 16'b1111111111111100;
		15'h3dd5: char_row_bitmap <= 16'b1111111111111100;
		15'h3dd6: char_row_bitmap <= 16'b1111111111111100;
		15'h3dd7: char_row_bitmap <= 16'b1111111111111100;
		15'h3dd8: char_row_bitmap <= 16'b1111111111111100;
		15'h3dd9: char_row_bitmap <= 16'b1111111111111100;
		15'h3dda: char_row_bitmap <= 16'b1111111111111100;
		15'h3ddb: char_row_bitmap <= 16'b1111111111111100;
		15'h3ddc: char_row_bitmap <= 16'b1111111111111100;
		15'h3ddd: char_row_bitmap <= 16'b1111111111111100;
		15'h3dde: char_row_bitmap <= 16'b1111111111111100;
		15'h3ddf: char_row_bitmap <= 16'b1111111111111100;
		15'h3de0: char_row_bitmap <= 16'b0000000000000000;
		15'h3de1: char_row_bitmap <= 16'b0000000000000000;
		15'h3de2: char_row_bitmap <= 16'b1111111111111100;
		15'h3de3: char_row_bitmap <= 16'b1111111111111100;
		15'h3de4: char_row_bitmap <= 16'b1111111111111100;
		15'h3de5: char_row_bitmap <= 16'b1111111111111100;
		15'h3de6: char_row_bitmap <= 16'b1111111111111100;
		15'h3de7: char_row_bitmap <= 16'b1111111111111100;
		15'h3de8: char_row_bitmap <= 16'b1111111111111100;
		15'h3de9: char_row_bitmap <= 16'b1111111111111100;
		15'h3dea: char_row_bitmap <= 16'b1111111111111100;
		15'h3deb: char_row_bitmap <= 16'b1111111111111100;
		15'h3dec: char_row_bitmap <= 16'b1111111111111100;
		15'h3ded: char_row_bitmap <= 16'b1111111111111100;
		15'h3dee: char_row_bitmap <= 16'b1111111111111100;
		15'h3def: char_row_bitmap <= 16'b1111111111111100;
		15'h3df0: char_row_bitmap <= 16'b1111111111111100;
		15'h3df1: char_row_bitmap <= 16'b1111111111111100;
		15'h3df2: char_row_bitmap <= 16'b1111111111111100;
		15'h3df3: char_row_bitmap <= 16'b1111111111111100;
		15'h3df4: char_row_bitmap <= 16'b1111111111111100;
		15'h3df5: char_row_bitmap <= 16'b1111111111111100;
		15'h3df6: char_row_bitmap <= 16'b1111111111111100;
		15'h3df7: char_row_bitmap <= 16'b1111111111111100;
		15'h3df8: char_row_bitmap <= 16'b1111111111111100;
		15'h3df9: char_row_bitmap <= 16'b1111111111111100;
		15'h3dfa: char_row_bitmap <= 16'b1111111111111100;
		15'h3dfb: char_row_bitmap <= 16'b1111111111111100;
		15'h3dfc: char_row_bitmap <= 16'b1111111111111100;
		15'h3dfd: char_row_bitmap <= 16'b1111111111111100;
		15'h3dfe: char_row_bitmap <= 16'b1111111111111100;
		15'h3dff: char_row_bitmap <= 16'b1111111111111100;
		15'h3e00: char_row_bitmap <= 16'b1111111111111100;
		15'h3e01: char_row_bitmap <= 16'b1111111111111100;
		15'h3e02: char_row_bitmap <= 16'b1111111111111100;
		15'h3e03: char_row_bitmap <= 16'b1111111111111100;
		15'h3e04: char_row_bitmap <= 16'b1111111111111100;
		15'h3e05: char_row_bitmap <= 16'b1111111111111100;
		15'h3e06: char_row_bitmap <= 16'b1111111111111100;
		15'h3e07: char_row_bitmap <= 16'b1111111111111100;
		15'h3e08: char_row_bitmap <= 16'b1111111111111111;
		15'h3e09: char_row_bitmap <= 16'b1111111111111111;
		15'h3e0a: char_row_bitmap <= 16'b0000000000000011;
		15'h3e0b: char_row_bitmap <= 16'b0000000000000011;
		15'h3e0c: char_row_bitmap <= 16'b0000000000000011;
		15'h3e0d: char_row_bitmap <= 16'b0000000000000011;
		15'h3e0e: char_row_bitmap <= 16'b0000000000000011;
		15'h3e0f: char_row_bitmap <= 16'b0000000000000011;
		15'h3e10: char_row_bitmap <= 16'b0000000000000011;
		15'h3e11: char_row_bitmap <= 16'b0000000000000011;
		15'h3e12: char_row_bitmap <= 16'b0000000000000011;
		15'h3e13: char_row_bitmap <= 16'b0000000000000011;
		15'h3e14: char_row_bitmap <= 16'b0000000000000011;
		15'h3e15: char_row_bitmap <= 16'b0000000000000011;
		15'h3e16: char_row_bitmap <= 16'b0000000000000011;
		15'h3e17: char_row_bitmap <= 16'b0000000000000011;
		15'h3e18: char_row_bitmap <= 16'b0000000000000011;
		15'h3e19: char_row_bitmap <= 16'b0000000000000011;
		15'h3e1a: char_row_bitmap <= 16'b1111111111111111;
		15'h3e1b: char_row_bitmap <= 16'b1111111111111111;
		15'h3e1c: char_row_bitmap <= 16'b1100000000000011;
		15'h3e1d: char_row_bitmap <= 16'b1100000000000011;
		15'h3e1e: char_row_bitmap <= 16'b1100000000000011;
		15'h3e1f: char_row_bitmap <= 16'b1100000000000011;
		15'h3e20: char_row_bitmap <= 16'b1100000000000011;
		15'h3e21: char_row_bitmap <= 16'b1100000000000011;
		15'h3e22: char_row_bitmap <= 16'b1100000000000011;
		15'h3e23: char_row_bitmap <= 16'b1100000000000011;
		15'h3e24: char_row_bitmap <= 16'b1100000000000011;
		15'h3e25: char_row_bitmap <= 16'b1100000000000011;
		15'h3e26: char_row_bitmap <= 16'b1100000000000011;
		15'h3e27: char_row_bitmap <= 16'b1100000000000011;
		15'h3e28: char_row_bitmap <= 16'b1100000000000011;
		15'h3e29: char_row_bitmap <= 16'b1100000000000011;
		15'h3e2a: char_row_bitmap <= 16'b1100000000000011;
		15'h3e2b: char_row_bitmap <= 16'b1100000000000011;
		15'h3e2c: char_row_bitmap <= 16'b1100000000000011;
		15'h3e2d: char_row_bitmap <= 16'b1100000000000011;
		15'h3e2e: char_row_bitmap <= 16'b1111111111111111;
		15'h3e2f: char_row_bitmap <= 16'b1111111111111111;
		15'h3e30: char_row_bitmap <= 16'b1111111111111111;
		15'h3e31: char_row_bitmap <= 16'b1111111111111111;
		15'h3e32: char_row_bitmap <= 16'b1100000000000000;
		15'h3e33: char_row_bitmap <= 16'b1100000000000000;
		15'h3e34: char_row_bitmap <= 16'b1100000000000000;
		15'h3e35: char_row_bitmap <= 16'b1100000000000000;
		15'h3e36: char_row_bitmap <= 16'b1100000000000000;
		15'h3e37: char_row_bitmap <= 16'b1100000000000000;
		15'h3e38: char_row_bitmap <= 16'b1100000000000000;
		15'h3e39: char_row_bitmap <= 16'b1100000000000000;
		15'h3e3a: char_row_bitmap <= 16'b1100000000000000;
		15'h3e3b: char_row_bitmap <= 16'b1100000000000000;
		15'h3e3c: char_row_bitmap <= 16'b1100000000000000;
		15'h3e3d: char_row_bitmap <= 16'b1100000000000000;
		15'h3e3e: char_row_bitmap <= 16'b1100000000000000;
		15'h3e3f: char_row_bitmap <= 16'b1100000000000000;
		15'h3e40: char_row_bitmap <= 16'b1100000000000000;
		15'h3e41: char_row_bitmap <= 16'b1100000000000000;
		15'h3e42: char_row_bitmap <= 16'b1111111111111111;
		15'h3e43: char_row_bitmap <= 16'b1111111111111111;
		15'h3e44: char_row_bitmap <= 16'b1111111111111111;
		15'h3e45: char_row_bitmap <= 16'b1111111111111111;
		15'h3e46: char_row_bitmap <= 16'b1100000000000011;
		15'h3e47: char_row_bitmap <= 16'b1100000000000011;
		15'h3e48: char_row_bitmap <= 16'b1100000000000011;
		15'h3e49: char_row_bitmap <= 16'b1100000000000011;
		15'h3e4a: char_row_bitmap <= 16'b1100000000000011;
		15'h3e4b: char_row_bitmap <= 16'b1100000000000011;
		15'h3e4c: char_row_bitmap <= 16'b1100000000000011;
		15'h3e4d: char_row_bitmap <= 16'b1100000000000011;
		15'h3e4e: char_row_bitmap <= 16'b1100000000000011;
		15'h3e4f: char_row_bitmap <= 16'b1100000000000011;
		15'h3e50: char_row_bitmap <= 16'b1100000000000011;
		15'h3e51: char_row_bitmap <= 16'b1100000000000011;
		15'h3e52: char_row_bitmap <= 16'b1100000000000011;
		15'h3e53: char_row_bitmap <= 16'b1100000000000011;
		15'h3e54: char_row_bitmap <= 16'b1100000000000011;
		15'h3e55: char_row_bitmap <= 16'b1100000000000011;
		15'h3e56: char_row_bitmap <= 16'b1100000000000011;
		15'h3e57: char_row_bitmap <= 16'b1100000000000011;
		15'h3e58: char_row_bitmap <= 16'b1111111111111111;
		15'h3e59: char_row_bitmap <= 16'b1111111111111111;
		15'h3e5a: char_row_bitmap <= 16'b1100000000000011;
		15'h3e5b: char_row_bitmap <= 16'b1100000000000011;
		15'h3e5c: char_row_bitmap <= 16'b1100000000000011;
		15'h3e5d: char_row_bitmap <= 16'b1100000000000011;
		15'h3e5e: char_row_bitmap <= 16'b1100000000000011;
		15'h3e5f: char_row_bitmap <= 16'b1100000000000011;
		15'h3e60: char_row_bitmap <= 16'b1100000000000011;
		15'h3e61: char_row_bitmap <= 16'b1100000000000011;
		15'h3e62: char_row_bitmap <= 16'b1100000000000011;
		15'h3e63: char_row_bitmap <= 16'b1100000000000011;
		15'h3e64: char_row_bitmap <= 16'b1100000000000011;
		15'h3e65: char_row_bitmap <= 16'b1100000000000011;
		15'h3e66: char_row_bitmap <= 16'b1100000000000011;
		15'h3e67: char_row_bitmap <= 16'b1100000000000011;
		15'h3e68: char_row_bitmap <= 16'b1100000000000011;
		15'h3e69: char_row_bitmap <= 16'b1100000000000011;
		15'h3e6a: char_row_bitmap <= 16'b1111111111111111;
		15'h3e6b: char_row_bitmap <= 16'b1111111111111111;
		15'h3e6c: char_row_bitmap <= 16'b0000000000000000;
		15'h3e6d: char_row_bitmap <= 16'b0000000000000000;
		15'h3e6e: char_row_bitmap <= 16'b0000000000000000;
		15'h3e6f: char_row_bitmap <= 16'b0000000000000000;
		15'h3e70: char_row_bitmap <= 16'b0000000000000000;
		15'h3e71: char_row_bitmap <= 16'b0000000000000000;
		15'h3e72: char_row_bitmap <= 16'b0000000000000000;
		15'h3e73: char_row_bitmap <= 16'b0000000000000000;
		15'h3e74: char_row_bitmap <= 16'b0000000000000000;
		15'h3e75: char_row_bitmap <= 16'b0000000000000000;
		15'h3e76: char_row_bitmap <= 16'b0000000000000000;
		15'h3e77: char_row_bitmap <= 16'b0000000000000000;
		15'h3e78: char_row_bitmap <= 16'b0000000000000000;
		15'h3e79: char_row_bitmap <= 16'b0000000000000000;
		15'h3e7a: char_row_bitmap <= 16'b0000000000000000;
		15'h3e7b: char_row_bitmap <= 16'b0000000000000000;
		15'h3e7c: char_row_bitmap <= 16'b0000000000000000;
		15'h3e7d: char_row_bitmap <= 16'b0000000000000000;
		15'h3e7e: char_row_bitmap <= 16'b0000000000000000;
		15'h3e7f: char_row_bitmap <= 16'b0000000000000000;
		15'h3e80: char_row_bitmap <= 16'b1111111111111111;
		15'h3e81: char_row_bitmap <= 16'b1111111111111111;
		15'h3e82: char_row_bitmap <= 16'b0000000000000000;
		15'h3e83: char_row_bitmap <= 16'b0000000000000000;
		15'h3e84: char_row_bitmap <= 16'b0000000000000000;
		15'h3e85: char_row_bitmap <= 16'b0000000000000000;
		15'h3e86: char_row_bitmap <= 16'b0000000000000000;
		15'h3e87: char_row_bitmap <= 16'b0000000000000000;
		15'h3e88: char_row_bitmap <= 16'b0000000000000000;
		15'h3e89: char_row_bitmap <= 16'b0000000000000000;
		15'h3e8a: char_row_bitmap <= 16'b0000000000000000;
		15'h3e8b: char_row_bitmap <= 16'b0000000000000000;
		15'h3e8c: char_row_bitmap <= 16'b0000000000000000;
		15'h3e8d: char_row_bitmap <= 16'b0000000000000000;
		15'h3e8e: char_row_bitmap <= 16'b0000000000000000;
		15'h3e8f: char_row_bitmap <= 16'b0000000000000000;
		15'h3e90: char_row_bitmap <= 16'b0000000000000000;
		15'h3e91: char_row_bitmap <= 16'b0000000000000000;
		15'h3e92: char_row_bitmap <= 16'b0000000000000000;
		15'h3e93: char_row_bitmap <= 16'b0000000000000000;
		15'h3e94: char_row_bitmap <= 16'b1111111111111111;
		15'h3e95: char_row_bitmap <= 16'b1111111111111111;
		15'h3e96: char_row_bitmap <= 16'b1111111111111111;
		15'h3e97: char_row_bitmap <= 16'b1111111111111111;
		15'h3e98: char_row_bitmap <= 16'b0000000000000000;
		15'h3e99: char_row_bitmap <= 16'b0000000000000000;
		15'h3e9a: char_row_bitmap <= 16'b0000000000000000;
		15'h3e9b: char_row_bitmap <= 16'b0000000000000000;
		15'h3e9c: char_row_bitmap <= 16'b0000000000000000;
		15'h3e9d: char_row_bitmap <= 16'b0000000000000000;
		15'h3e9e: char_row_bitmap <= 16'b0000000000000000;
		15'h3e9f: char_row_bitmap <= 16'b0000000000000000;
		15'h3ea0: char_row_bitmap <= 16'b0000000000000000;
		15'h3ea1: char_row_bitmap <= 16'b0000000000000000;
		15'h3ea2: char_row_bitmap <= 16'b0000000000000000;
		15'h3ea3: char_row_bitmap <= 16'b0000000000000000;
		15'h3ea4: char_row_bitmap <= 16'b0000000000000000;
		15'h3ea5: char_row_bitmap <= 16'b0000000000000000;
		15'h3ea6: char_row_bitmap <= 16'b0000000000000000;
		15'h3ea7: char_row_bitmap <= 16'b0000000000000000;
		15'h3ea8: char_row_bitmap <= 16'b1111111111111111;
		15'h3ea9: char_row_bitmap <= 16'b1111111111111111;
		15'h3eaa: char_row_bitmap <= 16'b1111111111111111;
		15'h3eab: char_row_bitmap <= 16'b1111111111111111;
		15'h3eac: char_row_bitmap <= 16'b1111111111111111;
		15'h3ead: char_row_bitmap <= 16'b1111111111111111;
		15'h3eae: char_row_bitmap <= 16'b0000000000000000;
		15'h3eaf: char_row_bitmap <= 16'b0000000000000000;
		15'h3eb0: char_row_bitmap <= 16'b0000000000000000;
		15'h3eb1: char_row_bitmap <= 16'b0000000000000000;
		15'h3eb2: char_row_bitmap <= 16'b0000000000000000;
		15'h3eb3: char_row_bitmap <= 16'b0000000000000000;
		15'h3eb4: char_row_bitmap <= 16'b0000000000000000;
		15'h3eb5: char_row_bitmap <= 16'b0000000000000000;
		15'h3eb6: char_row_bitmap <= 16'b0000000000000000;
		15'h3eb7: char_row_bitmap <= 16'b0000000000000000;
		15'h3eb8: char_row_bitmap <= 16'b0000000000000000;
		15'h3eb9: char_row_bitmap <= 16'b0000000000000000;
		15'h3eba: char_row_bitmap <= 16'b0000000000000000;
		15'h3ebb: char_row_bitmap <= 16'b0000000000000000;
		15'h3ebc: char_row_bitmap <= 16'b1111111111111111;
		15'h3ebd: char_row_bitmap <= 16'b1111111111111111;
		15'h3ebe: char_row_bitmap <= 16'b1111111111111111;
		15'h3ebf: char_row_bitmap <= 16'b1111111111111111;
		15'h3ec0: char_row_bitmap <= 16'b1111111111111111;
		15'h3ec1: char_row_bitmap <= 16'b1111111111111111;
		15'h3ec2: char_row_bitmap <= 16'b1111111111111111;
		15'h3ec3: char_row_bitmap <= 16'b1111111111111111;
		15'h3ec4: char_row_bitmap <= 16'b0000000000000000;
		15'h3ec5: char_row_bitmap <= 16'b0000000000000000;
		15'h3ec6: char_row_bitmap <= 16'b0000000000000000;
		15'h3ec7: char_row_bitmap <= 16'b0000000000000000;
		15'h3ec8: char_row_bitmap <= 16'b0000000000000000;
		15'h3ec9: char_row_bitmap <= 16'b0000000000000000;
		15'h3eca: char_row_bitmap <= 16'b0000000000000000;
		15'h3ecb: char_row_bitmap <= 16'b0000000000000000;
		15'h3ecc: char_row_bitmap <= 16'b0000000000000000;
		15'h3ecd: char_row_bitmap <= 16'b0000000000000000;
		15'h3ece: char_row_bitmap <= 16'b0000000000000000;
		15'h3ecf: char_row_bitmap <= 16'b0000000000000000;
		15'h3ed0: char_row_bitmap <= 16'b1111111111111111;
		15'h3ed1: char_row_bitmap <= 16'b1111111111111111;
		15'h3ed2: char_row_bitmap <= 16'b1111111111111111;
		15'h3ed3: char_row_bitmap <= 16'b1111111111111111;
		15'h3ed4: char_row_bitmap <= 16'b1111111111111111;
		15'h3ed5: char_row_bitmap <= 16'b1111111111111111;
		15'h3ed6: char_row_bitmap <= 16'b1111111111111111;
		15'h3ed7: char_row_bitmap <= 16'b1111111111111111;
		15'h3ed8: char_row_bitmap <= 16'b1111111111111111;
		15'h3ed9: char_row_bitmap <= 16'b1111111111111111;
		15'h3eda: char_row_bitmap <= 16'b0000000000000000;
		15'h3edb: char_row_bitmap <= 16'b0000000000000000;
		15'h3edc: char_row_bitmap <= 16'b0000000000000000;
		15'h3edd: char_row_bitmap <= 16'b0000000000000000;
		15'h3ede: char_row_bitmap <= 16'b0000000000000000;
		15'h3edf: char_row_bitmap <= 16'b0000000000000000;
		15'h3ee0: char_row_bitmap <= 16'b0000000000000000;
		15'h3ee1: char_row_bitmap <= 16'b0000000000000000;
		15'h3ee2: char_row_bitmap <= 16'b0000000000000000;
		15'h3ee3: char_row_bitmap <= 16'b0000000000000000;
		15'h3ee4: char_row_bitmap <= 16'b1111111111111111;
		15'h3ee5: char_row_bitmap <= 16'b1111111111111111;
		15'h3ee6: char_row_bitmap <= 16'b1111111111111111;
		15'h3ee7: char_row_bitmap <= 16'b1111111111111111;
		15'h3ee8: char_row_bitmap <= 16'b1111111111111111;
		15'h3ee9: char_row_bitmap <= 16'b1111111111111111;
		15'h3eea: char_row_bitmap <= 16'b1111111111111111;
		15'h3eeb: char_row_bitmap <= 16'b1111111111111111;
		15'h3eec: char_row_bitmap <= 16'b1111111111111111;
		15'h3eed: char_row_bitmap <= 16'b1111111111111111;
		15'h3eee: char_row_bitmap <= 16'b1111111111111111;
		15'h3eef: char_row_bitmap <= 16'b1111111111111111;
		15'h3ef0: char_row_bitmap <= 16'b0000000000000000;
		15'h3ef1: char_row_bitmap <= 16'b0000000000000000;
		15'h3ef2: char_row_bitmap <= 16'b0000000000000000;
		15'h3ef3: char_row_bitmap <= 16'b0000000000000000;
		15'h3ef4: char_row_bitmap <= 16'b0000000000000000;
		15'h3ef5: char_row_bitmap <= 16'b0000000000000000;
		15'h3ef6: char_row_bitmap <= 16'b0000000000000000;
		15'h3ef7: char_row_bitmap <= 16'b0000000000000000;
		15'h3ef8: char_row_bitmap <= 16'b1111111111111111;
		15'h3ef9: char_row_bitmap <= 16'b1111111111111111;
		15'h3efa: char_row_bitmap <= 16'b1111111111111111;
		15'h3efb: char_row_bitmap <= 16'b1111111111111111;
		15'h3efc: char_row_bitmap <= 16'b1111111111111111;
		15'h3efd: char_row_bitmap <= 16'b1111111111111111;
		15'h3efe: char_row_bitmap <= 16'b1111111111111111;
		15'h3eff: char_row_bitmap <= 16'b1111111111111111;
		15'h3f00: char_row_bitmap <= 16'b1111111111111111;
		15'h3f01: char_row_bitmap <= 16'b1111111111111111;
		15'h3f02: char_row_bitmap <= 16'b1111111111111111;
		15'h3f03: char_row_bitmap <= 16'b1111111111111111;
		15'h3f04: char_row_bitmap <= 16'b1111111111111111;
		15'h3f05: char_row_bitmap <= 16'b1111111111111111;
		15'h3f06: char_row_bitmap <= 16'b0000000000000000;
		15'h3f07: char_row_bitmap <= 16'b0000000000000000;
		15'h3f08: char_row_bitmap <= 16'b0000000000000000;
		15'h3f09: char_row_bitmap <= 16'b0000000000000000;
		15'h3f0a: char_row_bitmap <= 16'b0000000000000000;
		15'h3f0b: char_row_bitmap <= 16'b0000000000000000;
		15'h3f0c: char_row_bitmap <= 16'b1111111111111111;
		15'h3f0d: char_row_bitmap <= 16'b1111111111111111;
		15'h3f0e: char_row_bitmap <= 16'b1111111111111111;
		15'h3f0f: char_row_bitmap <= 16'b1111111111111111;
		15'h3f10: char_row_bitmap <= 16'b1111111111111111;
		15'h3f11: char_row_bitmap <= 16'b1111111111111111;
		15'h3f12: char_row_bitmap <= 16'b1111111111111111;
		15'h3f13: char_row_bitmap <= 16'b1111111111111111;
		15'h3f14: char_row_bitmap <= 16'b1111111111111111;
		15'h3f15: char_row_bitmap <= 16'b1111111111111111;
		15'h3f16: char_row_bitmap <= 16'b1111111111111111;
		15'h3f17: char_row_bitmap <= 16'b1111111111111111;
		15'h3f18: char_row_bitmap <= 16'b1111111111111111;
		15'h3f19: char_row_bitmap <= 16'b1111111111111111;
		15'h3f1a: char_row_bitmap <= 16'b1111111111111111;
		15'h3f1b: char_row_bitmap <= 16'b1111111111111111;
		15'h3f1c: char_row_bitmap <= 16'b0000000000000000;
		15'h3f1d: char_row_bitmap <= 16'b0000000000000000;
		15'h3f1e: char_row_bitmap <= 16'b0000000000000000;
		15'h3f1f: char_row_bitmap <= 16'b0000000000000000;
		15'h3f20: char_row_bitmap <= 16'b1111111111111111;
		15'h3f21: char_row_bitmap <= 16'b1111111111111111;
		15'h3f22: char_row_bitmap <= 16'b1111111111111111;
		15'h3f23: char_row_bitmap <= 16'b1111111111111111;
		15'h3f24: char_row_bitmap <= 16'b1111111111111111;
		15'h3f25: char_row_bitmap <= 16'b1111111111111111;
		15'h3f26: char_row_bitmap <= 16'b1111111111111111;
		15'h3f27: char_row_bitmap <= 16'b1111111111111111;
		15'h3f28: char_row_bitmap <= 16'b1111111111111111;
		15'h3f29: char_row_bitmap <= 16'b1111111111111111;
		15'h3f2a: char_row_bitmap <= 16'b1111111111111111;
		15'h3f2b: char_row_bitmap <= 16'b1111111111111111;
		15'h3f2c: char_row_bitmap <= 16'b1111111111111111;
		15'h3f2d: char_row_bitmap <= 16'b1111111111111111;
		15'h3f2e: char_row_bitmap <= 16'b1111111111111111;
		15'h3f2f: char_row_bitmap <= 16'b1111111111111111;
		15'h3f30: char_row_bitmap <= 16'b1111111111111111;
		15'h3f31: char_row_bitmap <= 16'b1111111111111111;
		15'h3f32: char_row_bitmap <= 16'b0000000000000000;
		15'h3f33: char_row_bitmap <= 16'b0000000000000000;
		15'h3f34: char_row_bitmap <= 16'b1111111111111111;
		15'h3f35: char_row_bitmap <= 16'b1111111111111111;
		15'h3f36: char_row_bitmap <= 16'b1111111111111111;
		15'h3f37: char_row_bitmap <= 16'b1111111111111111;
		15'h3f38: char_row_bitmap <= 16'b1111111111111111;
		15'h3f39: char_row_bitmap <= 16'b1111111111111111;
		15'h3f3a: char_row_bitmap <= 16'b1111111111111111;
		15'h3f3b: char_row_bitmap <= 16'b1111111111111111;
		15'h3f3c: char_row_bitmap <= 16'b1111111111111111;
		15'h3f3d: char_row_bitmap <= 16'b1111111111111111;
		15'h3f3e: char_row_bitmap <= 16'b1111111111111111;
		15'h3f3f: char_row_bitmap <= 16'b1111111111111111;
		15'h3f40: char_row_bitmap <= 16'b1111111111111111;
		15'h3f41: char_row_bitmap <= 16'b1111111111111111;
		15'h3f42: char_row_bitmap <= 16'b1111111111111111;
		15'h3f43: char_row_bitmap <= 16'b1111111111111111;
		15'h3f44: char_row_bitmap <= 16'b1111111111111111;
		15'h3f45: char_row_bitmap <= 16'b1111111111111111;
		15'h3f46: char_row_bitmap <= 16'b1111111111111111;
		15'h3f47: char_row_bitmap <= 16'b1111111111111111;
		15'h3f48: char_row_bitmap <= 16'b0000001111000000;
		15'h3f49: char_row_bitmap <= 16'b0000001111000000;
		15'h3f4a: char_row_bitmap <= 16'b0000001111000000;
		15'h3f4b: char_row_bitmap <= 16'b0000001111000000;
		15'h3f4c: char_row_bitmap <= 16'b0000011111100000;
		15'h3f4d: char_row_bitmap <= 16'b0001111111111000;
		15'h3f4e: char_row_bitmap <= 16'b0001110000111000;
		15'h3f4f: char_row_bitmap <= 16'b0011100000011100;
		15'h3f50: char_row_bitmap <= 16'b0011000000001100;
		15'h3f51: char_row_bitmap <= 16'b0011000000001100;
		15'h3f52: char_row_bitmap <= 16'b0011000000001100;
		15'h3f53: char_row_bitmap <= 16'b0011000000001100;
		15'h3f54: char_row_bitmap <= 16'b0011100000011100;
		15'h3f55: char_row_bitmap <= 16'b0001110000111000;
		15'h3f56: char_row_bitmap <= 16'b0001111111111000;
		15'h3f57: char_row_bitmap <= 16'b0000011111100000;
		15'h3f58: char_row_bitmap <= 16'b0000000000000000;
		15'h3f59: char_row_bitmap <= 16'b0000000000000000;
		15'h3f5a: char_row_bitmap <= 16'b0000000000000000;
		15'h3f5b: char_row_bitmap <= 16'b0000000000000000;
		15'h3f5c: char_row_bitmap <= 16'b0000000000000000;
		15'h3f5d: char_row_bitmap <= 16'b0000000000000000;
		15'h3f5e: char_row_bitmap <= 16'b0000000000000000;
		15'h3f5f: char_row_bitmap <= 16'b0000000000000000;
		15'h3f60: char_row_bitmap <= 16'b0000011111100000;
		15'h3f61: char_row_bitmap <= 16'b0001111111111000;
		15'h3f62: char_row_bitmap <= 16'b0001110000111000;
		15'h3f63: char_row_bitmap <= 16'b0011100000011100;
		15'h3f64: char_row_bitmap <= 16'b0011000000001111;
		15'h3f65: char_row_bitmap <= 16'b0011000000001111;
		15'h3f66: char_row_bitmap <= 16'b0011000000001111;
		15'h3f67: char_row_bitmap <= 16'b0011000000001111;
		15'h3f68: char_row_bitmap <= 16'b0011100000011100;
		15'h3f69: char_row_bitmap <= 16'b0001110000111000;
		15'h3f6a: char_row_bitmap <= 16'b0001111111111000;
		15'h3f6b: char_row_bitmap <= 16'b0000011111100000;
		15'h3f6c: char_row_bitmap <= 16'b0000000000000000;
		15'h3f6d: char_row_bitmap <= 16'b0000000000000000;
		15'h3f6e: char_row_bitmap <= 16'b0000000000000000;
		15'h3f6f: char_row_bitmap <= 16'b0000000000000000;
		15'h3f70: char_row_bitmap <= 16'b0000000000000000;
		15'h3f71: char_row_bitmap <= 16'b0000000000000000;
		15'h3f72: char_row_bitmap <= 16'b0000000000000000;
		15'h3f73: char_row_bitmap <= 16'b0000000000000000;
		15'h3f74: char_row_bitmap <= 16'b0000011111100000;
		15'h3f75: char_row_bitmap <= 16'b0001111111111000;
		15'h3f76: char_row_bitmap <= 16'b0001110000111000;
		15'h3f77: char_row_bitmap <= 16'b0011100000011100;
		15'h3f78: char_row_bitmap <= 16'b0011000000001100;
		15'h3f79: char_row_bitmap <= 16'b0011000000001100;
		15'h3f7a: char_row_bitmap <= 16'b0011000000001100;
		15'h3f7b: char_row_bitmap <= 16'b0011000000001100;
		15'h3f7c: char_row_bitmap <= 16'b0011100000011100;
		15'h3f7d: char_row_bitmap <= 16'b0001110000111000;
		15'h3f7e: char_row_bitmap <= 16'b0001111111111000;
		15'h3f7f: char_row_bitmap <= 16'b0000011111100000;
		15'h3f80: char_row_bitmap <= 16'b0000001111000000;
		15'h3f81: char_row_bitmap <= 16'b0000001111000000;
		15'h3f82: char_row_bitmap <= 16'b0000001111000000;
		15'h3f83: char_row_bitmap <= 16'b0000001111000000;
		15'h3f84: char_row_bitmap <= 16'b0000000000000000;
		15'h3f85: char_row_bitmap <= 16'b0000000000000000;
		15'h3f86: char_row_bitmap <= 16'b0000000000000000;
		15'h3f87: char_row_bitmap <= 16'b0000000000000000;
		15'h3f88: char_row_bitmap <= 16'b0000011111100000;
		15'h3f89: char_row_bitmap <= 16'b0001111111111000;
		15'h3f8a: char_row_bitmap <= 16'b0001110000111000;
		15'h3f8b: char_row_bitmap <= 16'b0011100000011100;
		15'h3f8c: char_row_bitmap <= 16'b1111000000001100;
		15'h3f8d: char_row_bitmap <= 16'b1111000000001100;
		15'h3f8e: char_row_bitmap <= 16'b1111000000001100;
		15'h3f8f: char_row_bitmap <= 16'b1111000000001100;
		15'h3f90: char_row_bitmap <= 16'b0011100000011100;
		15'h3f91: char_row_bitmap <= 16'b0001110000111000;
		15'h3f92: char_row_bitmap <= 16'b0001111111111000;
		15'h3f93: char_row_bitmap <= 16'b0000011111100000;
		15'h3f94: char_row_bitmap <= 16'b0000000000000000;
		15'h3f95: char_row_bitmap <= 16'b0000000000000000;
		15'h3f96: char_row_bitmap <= 16'b0000000000000000;
		15'h3f97: char_row_bitmap <= 16'b0000000000000000;
		15'h3f98: char_row_bitmap <= 16'b0000001111000000;
		15'h3f99: char_row_bitmap <= 16'b0000001111000000;
		15'h3f9a: char_row_bitmap <= 16'b0000001111000000;
		15'h3f9b: char_row_bitmap <= 16'b0000001111000000;
		15'h3f9c: char_row_bitmap <= 16'b0000011111100000;
		15'h3f9d: char_row_bitmap <= 16'b0001111111111000;
		15'h3f9e: char_row_bitmap <= 16'b0001110000111000;
		15'h3f9f: char_row_bitmap <= 16'b0011100000011100;
		15'h3fa0: char_row_bitmap <= 16'b0011000000001100;
		15'h3fa1: char_row_bitmap <= 16'b0011000000001100;
		15'h3fa2: char_row_bitmap <= 16'b0011000000001100;
		15'h3fa3: char_row_bitmap <= 16'b0011000000001100;
		15'h3fa4: char_row_bitmap <= 16'b0011100000011100;
		15'h3fa5: char_row_bitmap <= 16'b0001110000111000;
		15'h3fa6: char_row_bitmap <= 16'b0001111111111000;
		15'h3fa7: char_row_bitmap <= 16'b0000011111100000;
		15'h3fa8: char_row_bitmap <= 16'b0000001111000000;
		15'h3fa9: char_row_bitmap <= 16'b0000001111000000;
		15'h3faa: char_row_bitmap <= 16'b0000001111000000;
		15'h3fab: char_row_bitmap <= 16'b0000001111000000;
		15'h3fac: char_row_bitmap <= 16'b0000000000000000;
		15'h3fad: char_row_bitmap <= 16'b0000000000000000;
		15'h3fae: char_row_bitmap <= 16'b0000000000000000;
		15'h3faf: char_row_bitmap <= 16'b0000000000000000;
		15'h3fb0: char_row_bitmap <= 16'b0000011111100000;
		15'h3fb1: char_row_bitmap <= 16'b0001111111111000;
		15'h3fb2: char_row_bitmap <= 16'b0001110000111000;
		15'h3fb3: char_row_bitmap <= 16'b0011100000011100;
		15'h3fb4: char_row_bitmap <= 16'b1111000000001111;
		15'h3fb5: char_row_bitmap <= 16'b1111000000001111;
		15'h3fb6: char_row_bitmap <= 16'b1111000000001111;
		15'h3fb7: char_row_bitmap <= 16'b1111000000001111;
		15'h3fb8: char_row_bitmap <= 16'b0011100000011100;
		15'h3fb9: char_row_bitmap <= 16'b0001110000111000;
		15'h3fba: char_row_bitmap <= 16'b0001111111111000;
		15'h3fbb: char_row_bitmap <= 16'b0000011111100000;
		15'h3fbc: char_row_bitmap <= 16'b0000000000000000;
		15'h3fbd: char_row_bitmap <= 16'b0000000000000000;
		15'h3fbe: char_row_bitmap <= 16'b0000000000000000;
		15'h3fbf: char_row_bitmap <= 16'b0000000000000000;
		15'h3fc0: char_row_bitmap <= 16'b1111111111111100;
		15'h3fc1: char_row_bitmap <= 16'b1111111111111100;
		15'h3fc2: char_row_bitmap <= 16'b0000000000000000;
		15'h3fc3: char_row_bitmap <= 16'b0000000000000000;
		15'h3fc4: char_row_bitmap <= 16'b0000000000000000;
		15'h3fc5: char_row_bitmap <= 16'b0000000000000000;
		15'h3fc6: char_row_bitmap <= 16'b0000000000000000;
		15'h3fc7: char_row_bitmap <= 16'b0000000000000000;
		15'h3fc8: char_row_bitmap <= 16'b0000000000000000;
		15'h3fc9: char_row_bitmap <= 16'b0000000000000000;
		15'h3fca: char_row_bitmap <= 16'b0000000000000000;
		15'h3fcb: char_row_bitmap <= 16'b0000000000000000;
		15'h3fcc: char_row_bitmap <= 16'b0000000000000000;
		15'h3fcd: char_row_bitmap <= 16'b0000000000000000;
		15'h3fce: char_row_bitmap <= 16'b0000000000000000;
		15'h3fcf: char_row_bitmap <= 16'b0000000000000000;
		15'h3fd0: char_row_bitmap <= 16'b0000000000000000;
		15'h3fd1: char_row_bitmap <= 16'b0000000000000000;
		15'h3fd2: char_row_bitmap <= 16'b0000000000000000;
		15'h3fd3: char_row_bitmap <= 16'b0000000000000000;
		15'h3fd4: char_row_bitmap <= 16'b1111111111111100;
		15'h3fd5: char_row_bitmap <= 16'b1111111111111100;
		15'h3fd6: char_row_bitmap <= 16'b1111111111111100;
		15'h3fd7: char_row_bitmap <= 16'b1111111111111100;
		15'h3fd8: char_row_bitmap <= 16'b0000000000000000;
		15'h3fd9: char_row_bitmap <= 16'b0000000000000000;
		15'h3fda: char_row_bitmap <= 16'b0000000000000000;
		15'h3fdb: char_row_bitmap <= 16'b0000000000000000;
		15'h3fdc: char_row_bitmap <= 16'b0000000000000000;
		15'h3fdd: char_row_bitmap <= 16'b0000000000000000;
		15'h3fde: char_row_bitmap <= 16'b0000000000000000;
		15'h3fdf: char_row_bitmap <= 16'b0000000000000000;
		15'h3fe0: char_row_bitmap <= 16'b0000000000000000;
		15'h3fe1: char_row_bitmap <= 16'b0000000000000000;
		15'h3fe2: char_row_bitmap <= 16'b0000000000000000;
		15'h3fe3: char_row_bitmap <= 16'b0000000000000000;
		15'h3fe4: char_row_bitmap <= 16'b0000000000000000;
		15'h3fe5: char_row_bitmap <= 16'b0000000000000000;
		15'h3fe6: char_row_bitmap <= 16'b0000000000000000;
		15'h3fe7: char_row_bitmap <= 16'b0000000000000000;
		15'h3fe8: char_row_bitmap <= 16'b1111111111111100;
		15'h3fe9: char_row_bitmap <= 16'b1111111111111100;
		15'h3fea: char_row_bitmap <= 16'b1111111111111100;
		15'h3feb: char_row_bitmap <= 16'b1111111111111100;
		15'h3fec: char_row_bitmap <= 16'b1111111111111100;
		15'h3fed: char_row_bitmap <= 16'b1111111111111100;
		15'h3fee: char_row_bitmap <= 16'b0000000000000000;
		15'h3fef: char_row_bitmap <= 16'b0000000000000000;
		15'h3ff0: char_row_bitmap <= 16'b0000000000000000;
		15'h3ff1: char_row_bitmap <= 16'b0000000000000000;
		15'h3ff2: char_row_bitmap <= 16'b0000000000000000;
		15'h3ff3: char_row_bitmap <= 16'b0000000000000000;
		15'h3ff4: char_row_bitmap <= 16'b0000000000000000;
		15'h3ff5: char_row_bitmap <= 16'b0000000000000000;
		15'h3ff6: char_row_bitmap <= 16'b0000000000000000;
		15'h3ff7: char_row_bitmap <= 16'b0000000000000000;
		15'h3ff8: char_row_bitmap <= 16'b0000000000000000;
		15'h3ff9: char_row_bitmap <= 16'b0000000000000000;
		15'h3ffa: char_row_bitmap <= 16'b0000000000000000;
		15'h3ffb: char_row_bitmap <= 16'b0000000000000000;
		15'h3ffc: char_row_bitmap <= 16'b1111111111111100;
		15'h3ffd: char_row_bitmap <= 16'b1111111111111100;
		15'h3ffe: char_row_bitmap <= 16'b1111111111111100;
		15'h3fff: char_row_bitmap <= 16'b1111111111111100;
		15'h4000: char_row_bitmap <= 16'b1111111111111100;
		15'h4001: char_row_bitmap <= 16'b1111111111111100;
		15'h4002: char_row_bitmap <= 16'b1111111111111100;
		15'h4003: char_row_bitmap <= 16'b1111111111111100;
		15'h4004: char_row_bitmap <= 16'b0000000000000000;
		15'h4005: char_row_bitmap <= 16'b0000000000000000;
		15'h4006: char_row_bitmap <= 16'b0000000000000000;
		15'h4007: char_row_bitmap <= 16'b0000000000000000;
		15'h4008: char_row_bitmap <= 16'b0000000000000000;
		15'h4009: char_row_bitmap <= 16'b0000000000000000;
		15'h400a: char_row_bitmap <= 16'b0000000000000000;
		15'h400b: char_row_bitmap <= 16'b0000000000000000;
		15'h400c: char_row_bitmap <= 16'b0000000000000000;
		15'h400d: char_row_bitmap <= 16'b0000000000000000;
		15'h400e: char_row_bitmap <= 16'b0000000000000000;
		15'h400f: char_row_bitmap <= 16'b0000000000000000;
		15'h4010: char_row_bitmap <= 16'b1111111111111100;
		15'h4011: char_row_bitmap <= 16'b1111111111111100;
		15'h4012: char_row_bitmap <= 16'b1111111111111100;
		15'h4013: char_row_bitmap <= 16'b1111111111111100;
		15'h4014: char_row_bitmap <= 16'b1111111111111100;
		15'h4015: char_row_bitmap <= 16'b1111111111111100;
		15'h4016: char_row_bitmap <= 16'b1111111111111100;
		15'h4017: char_row_bitmap <= 16'b1111111111111100;
		15'h4018: char_row_bitmap <= 16'b1111111111111100;
		15'h4019: char_row_bitmap <= 16'b1111111111111100;
		15'h401a: char_row_bitmap <= 16'b0000000000000000;
		15'h401b: char_row_bitmap <= 16'b0000000000000000;
		15'h401c: char_row_bitmap <= 16'b0000000000000000;
		15'h401d: char_row_bitmap <= 16'b0000000000000000;
		15'h401e: char_row_bitmap <= 16'b0000000000000000;
		15'h401f: char_row_bitmap <= 16'b0000000000000000;
		15'h4020: char_row_bitmap <= 16'b0000000000000000;
		15'h4021: char_row_bitmap <= 16'b0000000000000000;
		15'h4022: char_row_bitmap <= 16'b0000000000000000;
		15'h4023: char_row_bitmap <= 16'b0000000000000000;
		15'h4024: char_row_bitmap <= 16'b1111111111111100;
		15'h4025: char_row_bitmap <= 16'b1111111111111100;
		15'h4026: char_row_bitmap <= 16'b1111111111111100;
		15'h4027: char_row_bitmap <= 16'b1111111111111100;
		15'h4028: char_row_bitmap <= 16'b1111111111111100;
		15'h4029: char_row_bitmap <= 16'b1111111111111100;
		15'h402a: char_row_bitmap <= 16'b1111111111111100;
		15'h402b: char_row_bitmap <= 16'b1111111111111100;
		15'h402c: char_row_bitmap <= 16'b1111111111111100;
		15'h402d: char_row_bitmap <= 16'b1111111111111100;
		15'h402e: char_row_bitmap <= 16'b1111111111111100;
		15'h402f: char_row_bitmap <= 16'b1111111111111100;
		15'h4030: char_row_bitmap <= 16'b0000000000000000;
		15'h4031: char_row_bitmap <= 16'b0000000000000000;
		15'h4032: char_row_bitmap <= 16'b0000000000000000;
		15'h4033: char_row_bitmap <= 16'b0000000000000000;
		15'h4034: char_row_bitmap <= 16'b0000000000000000;
		15'h4035: char_row_bitmap <= 16'b0000000000000000;
		15'h4036: char_row_bitmap <= 16'b0000000000000000;
		15'h4037: char_row_bitmap <= 16'b0000000000000000;
		15'h4038: char_row_bitmap <= 16'b1111111111111100;
		15'h4039: char_row_bitmap <= 16'b1111111111111100;
		15'h403a: char_row_bitmap <= 16'b1111111111111100;
		15'h403b: char_row_bitmap <= 16'b1111111111111100;
		15'h403c: char_row_bitmap <= 16'b1111111111111100;
		15'h403d: char_row_bitmap <= 16'b1111111111111100;
		15'h403e: char_row_bitmap <= 16'b1111111111111100;
		15'h403f: char_row_bitmap <= 16'b1111111111111100;
		15'h4040: char_row_bitmap <= 16'b1111111111111100;
		15'h4041: char_row_bitmap <= 16'b1111111111111100;
		15'h4042: char_row_bitmap <= 16'b1111111111111100;
		15'h4043: char_row_bitmap <= 16'b1111111111111100;
		15'h4044: char_row_bitmap <= 16'b1111111111111100;
		15'h4045: char_row_bitmap <= 16'b1111111111111100;
		15'h4046: char_row_bitmap <= 16'b0000000000000000;
		15'h4047: char_row_bitmap <= 16'b0000000000000000;
		15'h4048: char_row_bitmap <= 16'b0000000000000000;
		15'h4049: char_row_bitmap <= 16'b0000000000000000;
		15'h404a: char_row_bitmap <= 16'b0000000000000000;
		15'h404b: char_row_bitmap <= 16'b0000000000000000;
		15'h404c: char_row_bitmap <= 16'b1111111111111100;
		15'h404d: char_row_bitmap <= 16'b1111111111111100;
		15'h404e: char_row_bitmap <= 16'b1111111111111100;
		15'h404f: char_row_bitmap <= 16'b1111111111111100;
		15'h4050: char_row_bitmap <= 16'b1111111111111100;
		15'h4051: char_row_bitmap <= 16'b1111111111111100;
		15'h4052: char_row_bitmap <= 16'b1111111111111100;
		15'h4053: char_row_bitmap <= 16'b1111111111111100;
		15'h4054: char_row_bitmap <= 16'b1111111111111100;
		15'h4055: char_row_bitmap <= 16'b1111111111111100;
		15'h4056: char_row_bitmap <= 16'b1111111111111100;
		15'h4057: char_row_bitmap <= 16'b1111111111111100;
		15'h4058: char_row_bitmap <= 16'b1111111111111100;
		15'h4059: char_row_bitmap <= 16'b1111111111111100;
		15'h405a: char_row_bitmap <= 16'b1111111111111100;
		15'h405b: char_row_bitmap <= 16'b1111111111111100;
		15'h405c: char_row_bitmap <= 16'b0000000000000000;
		15'h405d: char_row_bitmap <= 16'b0000000000000000;
		15'h405e: char_row_bitmap <= 16'b0000000000000000;
		15'h405f: char_row_bitmap <= 16'b0000000000000000;
		15'h4060: char_row_bitmap <= 16'b1111111111111100;
		15'h4061: char_row_bitmap <= 16'b1111111111111100;
		15'h4062: char_row_bitmap <= 16'b1111111111111100;
		15'h4063: char_row_bitmap <= 16'b1111111111111100;
		15'h4064: char_row_bitmap <= 16'b1111111111111100;
		15'h4065: char_row_bitmap <= 16'b1111111111111100;
		15'h4066: char_row_bitmap <= 16'b1111111111111100;
		15'h4067: char_row_bitmap <= 16'b1111111111111100;
		15'h4068: char_row_bitmap <= 16'b1111111111111100;
		15'h4069: char_row_bitmap <= 16'b1111111111111100;
		15'h406a: char_row_bitmap <= 16'b1111111111111100;
		15'h406b: char_row_bitmap <= 16'b1111111111111100;
		15'h406c: char_row_bitmap <= 16'b1111111111111100;
		15'h406d: char_row_bitmap <= 16'b1111111111111100;
		15'h406e: char_row_bitmap <= 16'b1111111111111100;
		15'h406f: char_row_bitmap <= 16'b1111111111111100;
		15'h4070: char_row_bitmap <= 16'b1111111111111100;
		15'h4071: char_row_bitmap <= 16'b1111111111111100;
		15'h4072: char_row_bitmap <= 16'b0000000000000000;
		15'h4073: char_row_bitmap <= 16'b0000000000000000;
		15'h4074: char_row_bitmap <= 16'b1111111111111100;
		15'h4075: char_row_bitmap <= 16'b1111111111111100;
		15'h4076: char_row_bitmap <= 16'b1111111111111100;
		15'h4077: char_row_bitmap <= 16'b1111111111111100;
		15'h4078: char_row_bitmap <= 16'b1111111111111100;
		15'h4079: char_row_bitmap <= 16'b1111111111111100;
		15'h407a: char_row_bitmap <= 16'b1111111111111100;
		15'h407b: char_row_bitmap <= 16'b1111111111111100;
		15'h407c: char_row_bitmap <= 16'b1111111111111100;
		15'h407d: char_row_bitmap <= 16'b1111111111111100;
		15'h407e: char_row_bitmap <= 16'b1111111111111100;
		15'h407f: char_row_bitmap <= 16'b1111111111111100;
		15'h4080: char_row_bitmap <= 16'b1111111111111100;
		15'h4081: char_row_bitmap <= 16'b1111111111111100;
		15'h4082: char_row_bitmap <= 16'b1111111111111100;
		15'h4083: char_row_bitmap <= 16'b1111111111111100;
		15'h4084: char_row_bitmap <= 16'b1111111111111100;
		15'h4085: char_row_bitmap <= 16'b1111111111111100;
		15'h4086: char_row_bitmap <= 16'b1111111111111100;
		15'h4087: char_row_bitmap <= 16'b1111111111111100;
		15'h4088: char_row_bitmap <= 16'b0000001111000000;
		15'h4089: char_row_bitmap <= 16'b0000001111000000;
		15'h408a: char_row_bitmap <= 16'b0000001111000000;
		15'h408b: char_row_bitmap <= 16'b0000001111000000;
		15'h408c: char_row_bitmap <= 16'b0000011111100000;
		15'h408d: char_row_bitmap <= 16'b0001111111111000;
		15'h408e: char_row_bitmap <= 16'b0001111111111000;
		15'h408f: char_row_bitmap <= 16'b0011111111111100;
		15'h4090: char_row_bitmap <= 16'b0011111111111100;
		15'h4091: char_row_bitmap <= 16'b0011111111111100;
		15'h4092: char_row_bitmap <= 16'b0011111111111100;
		15'h4093: char_row_bitmap <= 16'b0011111111111100;
		15'h4094: char_row_bitmap <= 16'b0011111111111100;
		15'h4095: char_row_bitmap <= 16'b0001111111111000;
		15'h4096: char_row_bitmap <= 16'b0001111111111000;
		15'h4097: char_row_bitmap <= 16'b0000011111100000;
		15'h4098: char_row_bitmap <= 16'b0000000000000000;
		15'h4099: char_row_bitmap <= 16'b0000000000000000;
		15'h409a: char_row_bitmap <= 16'b0000000000000000;
		15'h409b: char_row_bitmap <= 16'b0000000000000000;
		15'h409c: char_row_bitmap <= 16'b0000000000000000;
		15'h409d: char_row_bitmap <= 16'b0000000000000000;
		15'h409e: char_row_bitmap <= 16'b0000000000000000;
		15'h409f: char_row_bitmap <= 16'b0000000000000000;
		15'h40a0: char_row_bitmap <= 16'b0000011111100000;
		15'h40a1: char_row_bitmap <= 16'b0001111111111000;
		15'h40a2: char_row_bitmap <= 16'b0001111111111000;
		15'h40a3: char_row_bitmap <= 16'b0011111111111100;
		15'h40a4: char_row_bitmap <= 16'b0011111111111111;
		15'h40a5: char_row_bitmap <= 16'b0011111111111111;
		15'h40a6: char_row_bitmap <= 16'b0011111111111111;
		15'h40a7: char_row_bitmap <= 16'b0011111111111111;
		15'h40a8: char_row_bitmap <= 16'b0011111111111100;
		15'h40a9: char_row_bitmap <= 16'b0001111111111000;
		15'h40aa: char_row_bitmap <= 16'b0001111111111000;
		15'h40ab: char_row_bitmap <= 16'b0000011111100000;
		15'h40ac: char_row_bitmap <= 16'b0000000000000000;
		15'h40ad: char_row_bitmap <= 16'b0000000000000000;
		15'h40ae: char_row_bitmap <= 16'b0000000000000000;
		15'h40af: char_row_bitmap <= 16'b0000000000000000;
		15'h40b0: char_row_bitmap <= 16'b0000000000000000;
		15'h40b1: char_row_bitmap <= 16'b0000000000000000;
		15'h40b2: char_row_bitmap <= 16'b0000000000000000;
		15'h40b3: char_row_bitmap <= 16'b0000000000000000;
		15'h40b4: char_row_bitmap <= 16'b0000011111100000;
		15'h40b5: char_row_bitmap <= 16'b0001111111111000;
		15'h40b6: char_row_bitmap <= 16'b0001111111111000;
		15'h40b7: char_row_bitmap <= 16'b0011111111111100;
		15'h40b8: char_row_bitmap <= 16'b0011111111111100;
		15'h40b9: char_row_bitmap <= 16'b0011111111111100;
		15'h40ba: char_row_bitmap <= 16'b0011111111111100;
		15'h40bb: char_row_bitmap <= 16'b0011111111111100;
		15'h40bc: char_row_bitmap <= 16'b0011111111111100;
		15'h40bd: char_row_bitmap <= 16'b0001111111111000;
		15'h40be: char_row_bitmap <= 16'b0001111111111000;
		15'h40bf: char_row_bitmap <= 16'b0000011111100000;
		15'h40c0: char_row_bitmap <= 16'b0000001111000000;
		15'h40c1: char_row_bitmap <= 16'b0000001111000000;
		15'h40c2: char_row_bitmap <= 16'b0000001111000000;
		15'h40c3: char_row_bitmap <= 16'b0000001111000000;
		15'h40c4: char_row_bitmap <= 16'b0000000000000000;
		15'h40c5: char_row_bitmap <= 16'b0000000000000000;
		15'h40c6: char_row_bitmap <= 16'b0000000000000000;
		15'h40c7: char_row_bitmap <= 16'b0000000000000000;
		15'h40c8: char_row_bitmap <= 16'b0000011111100000;
		15'h40c9: char_row_bitmap <= 16'b0001111111111000;
		15'h40ca: char_row_bitmap <= 16'b0001111111111000;
		15'h40cb: char_row_bitmap <= 16'b0011111111111100;
		15'h40cc: char_row_bitmap <= 16'b1111111111111100;
		15'h40cd: char_row_bitmap <= 16'b1111111111111100;
		15'h40ce: char_row_bitmap <= 16'b1111111111111100;
		15'h40cf: char_row_bitmap <= 16'b1111111111111100;
		15'h40d0: char_row_bitmap <= 16'b0011111111111100;
		15'h40d1: char_row_bitmap <= 16'b0001111111111000;
		15'h40d2: char_row_bitmap <= 16'b0001111111111000;
		15'h40d3: char_row_bitmap <= 16'b0000011111100000;
		15'h40d4: char_row_bitmap <= 16'b0000000000000000;
		15'h40d5: char_row_bitmap <= 16'b0000000000000000;
		15'h40d6: char_row_bitmap <= 16'b0000000000000000;
		15'h40d7: char_row_bitmap <= 16'b0000000000000000;
		15'h40d8: char_row_bitmap <= 16'b0000001111000000;
		15'h40d9: char_row_bitmap <= 16'b0000001111000000;
		15'h40da: char_row_bitmap <= 16'b0000001111000000;
		15'h40db: char_row_bitmap <= 16'b0000001111000000;
		15'h40dc: char_row_bitmap <= 16'b0000011111100000;
		15'h40dd: char_row_bitmap <= 16'b0001111111111000;
		15'h40de: char_row_bitmap <= 16'b0001111111111000;
		15'h40df: char_row_bitmap <= 16'b0011111111111100;
		15'h40e0: char_row_bitmap <= 16'b0011111111111100;
		15'h40e1: char_row_bitmap <= 16'b0011111111111100;
		15'h40e2: char_row_bitmap <= 16'b0011111111111100;
		15'h40e3: char_row_bitmap <= 16'b0011111111111100;
		15'h40e4: char_row_bitmap <= 16'b0011111111111100;
		15'h40e5: char_row_bitmap <= 16'b0001111111111000;
		15'h40e6: char_row_bitmap <= 16'b0001111111111000;
		15'h40e7: char_row_bitmap <= 16'b0000011111100000;
		15'h40e8: char_row_bitmap <= 16'b0000001111000000;
		15'h40e9: char_row_bitmap <= 16'b0000001111000000;
		15'h40ea: char_row_bitmap <= 16'b0000001111000000;
		15'h40eb: char_row_bitmap <= 16'b0000001111000000;
		15'h40ec: char_row_bitmap <= 16'b0000000000000000;
		15'h40ed: char_row_bitmap <= 16'b0000000000000000;
		15'h40ee: char_row_bitmap <= 16'b0000000000000000;
		15'h40ef: char_row_bitmap <= 16'b0000000000000000;
		15'h40f0: char_row_bitmap <= 16'b0000011111100000;
		15'h40f1: char_row_bitmap <= 16'b0001111111111000;
		15'h40f2: char_row_bitmap <= 16'b0001111111111000;
		15'h40f3: char_row_bitmap <= 16'b0011111111111100;
		15'h40f4: char_row_bitmap <= 16'b1111111111111111;
		15'h40f5: char_row_bitmap <= 16'b1111111111111111;
		15'h40f6: char_row_bitmap <= 16'b1111111111111111;
		15'h40f7: char_row_bitmap <= 16'b1111111111111111;
		15'h40f8: char_row_bitmap <= 16'b0011111111111100;
		15'h40f9: char_row_bitmap <= 16'b0001111111111000;
		15'h40fa: char_row_bitmap <= 16'b0001111111111000;
		15'h40fb: char_row_bitmap <= 16'b0000011111100000;
		15'h40fc: char_row_bitmap <= 16'b0000000000000000;
		15'h40fd: char_row_bitmap <= 16'b0000000000000000;
		15'h40fe: char_row_bitmap <= 16'b0000000000000000;
		15'h40ff: char_row_bitmap <= 16'b0000000000000000;
		15'h4100: char_row_bitmap <= 16'b0000000000000000;
		15'h4101: char_row_bitmap <= 16'b0000000000000000;
		15'h4102: char_row_bitmap <= 16'b0000001111000000;
		15'h4103: char_row_bitmap <= 16'b0000111111110000;
		15'h4104: char_row_bitmap <= 16'b0001111111111000;
		15'h4105: char_row_bitmap <= 16'b0001111111111000;
		15'h4106: char_row_bitmap <= 16'b0011111111111100;
		15'h4107: char_row_bitmap <= 16'b0011111111111100;
		15'h4108: char_row_bitmap <= 16'b0111111111111110;
		15'h4109: char_row_bitmap <= 16'b0111111111111110;
		15'h410a: char_row_bitmap <= 16'b0111111111111110;
		15'h410b: char_row_bitmap <= 16'b0111111111111110;
		15'h410c: char_row_bitmap <= 16'b0111111111111110;
		15'h410d: char_row_bitmap <= 16'b1111111111111111;
		15'h410e: char_row_bitmap <= 16'b1111111111111111;
		15'h410f: char_row_bitmap <= 16'b1111111111111111;
		15'h4110: char_row_bitmap <= 16'b1111111111111111;
		15'h4111: char_row_bitmap <= 16'b1111111111111111;
		15'h4112: char_row_bitmap <= 16'b1111111111111111;
		15'h4113: char_row_bitmap <= 16'b1111111111111111;
		15'h4114: char_row_bitmap <= 16'b1111000000000000;
		15'h4115: char_row_bitmap <= 16'b1111111100000000;
		15'h4116: char_row_bitmap <= 16'b1111111111000000;
		15'h4117: char_row_bitmap <= 16'b1111111111110000;
		15'h4118: char_row_bitmap <= 16'b1111111111111000;
		15'h4119: char_row_bitmap <= 16'b1111111111111000;
		15'h411a: char_row_bitmap <= 16'b1111111111111100;
		15'h411b: char_row_bitmap <= 16'b1111111111111100;
		15'h411c: char_row_bitmap <= 16'b1111111111111110;
		15'h411d: char_row_bitmap <= 16'b1111111111111110;
		15'h411e: char_row_bitmap <= 16'b1111111111111110;
		15'h411f: char_row_bitmap <= 16'b1111111111111110;
		15'h4120: char_row_bitmap <= 16'b1111111111111100;
		15'h4121: char_row_bitmap <= 16'b1111111111111100;
		15'h4122: char_row_bitmap <= 16'b1111111111111000;
		15'h4123: char_row_bitmap <= 16'b1111111111111000;
		15'h4124: char_row_bitmap <= 16'b1111111111110000;
		15'h4125: char_row_bitmap <= 16'b1111111111000000;
		15'h4126: char_row_bitmap <= 16'b1111111100000000;
		15'h4127: char_row_bitmap <= 16'b1111000000000000;
		15'h4128: char_row_bitmap <= 16'b1111111111111111;
		15'h4129: char_row_bitmap <= 16'b1111111111111111;
		15'h412a: char_row_bitmap <= 16'b1111111111111111;
		15'h412b: char_row_bitmap <= 16'b1111111111111111;
		15'h412c: char_row_bitmap <= 16'b1111111111111111;
		15'h412d: char_row_bitmap <= 16'b1111111111111111;
		15'h412e: char_row_bitmap <= 16'b1111111111111111;
		15'h412f: char_row_bitmap <= 16'b0111111111111110;
		15'h4130: char_row_bitmap <= 16'b0111111111111110;
		15'h4131: char_row_bitmap <= 16'b0111111111111110;
		15'h4132: char_row_bitmap <= 16'b0111111111111110;
		15'h4133: char_row_bitmap <= 16'b0111111111111110;
		15'h4134: char_row_bitmap <= 16'b0011111111111100;
		15'h4135: char_row_bitmap <= 16'b0011111111111100;
		15'h4136: char_row_bitmap <= 16'b0001111111111000;
		15'h4137: char_row_bitmap <= 16'b0001111111111000;
		15'h4138: char_row_bitmap <= 16'b0000111111110000;
		15'h4139: char_row_bitmap <= 16'b0000001111000000;
		15'h413a: char_row_bitmap <= 16'b0000000000000000;
		15'h413b: char_row_bitmap <= 16'b0000000000000000;
		15'h413c: char_row_bitmap <= 16'b0000000000001111;
		15'h413d: char_row_bitmap <= 16'b0000000011111111;
		15'h413e: char_row_bitmap <= 16'b0000001111111111;
		15'h413f: char_row_bitmap <= 16'b0000111111111111;
		15'h4140: char_row_bitmap <= 16'b0001111111111111;
		15'h4141: char_row_bitmap <= 16'b0001111111111111;
		15'h4142: char_row_bitmap <= 16'b0011111111111111;
		15'h4143: char_row_bitmap <= 16'b0011111111111111;
		15'h4144: char_row_bitmap <= 16'b0111111111111111;
		15'h4145: char_row_bitmap <= 16'b0111111111111111;
		15'h4146: char_row_bitmap <= 16'b0111111111111111;
		15'h4147: char_row_bitmap <= 16'b0111111111111111;
		15'h4148: char_row_bitmap <= 16'b0011111111111111;
		15'h4149: char_row_bitmap <= 16'b0011111111111111;
		15'h414a: char_row_bitmap <= 16'b0001111111111111;
		15'h414b: char_row_bitmap <= 16'b0001111111111111;
		15'h414c: char_row_bitmap <= 16'b0000111111111111;
		15'h414d: char_row_bitmap <= 16'b0000001111111111;
		15'h414e: char_row_bitmap <= 16'b0000000011111111;
		15'h414f: char_row_bitmap <= 16'b0000000000001111;
		15'h4150: char_row_bitmap <= 16'b1111000000000000;
		15'h4151: char_row_bitmap <= 16'b1111111100000000;
		15'h4152: char_row_bitmap <= 16'b1111111111000000;
		15'h4153: char_row_bitmap <= 16'b1111111111100000;
		15'h4154: char_row_bitmap <= 16'b1111111111110000;
		15'h4155: char_row_bitmap <= 16'b1111111111111000;
		15'h4156: char_row_bitmap <= 16'b1111111111111100;
		15'h4157: char_row_bitmap <= 16'b1111111111111100;
		15'h4158: char_row_bitmap <= 16'b1111111111111100;
		15'h4159: char_row_bitmap <= 16'b1111111111111110;
		15'h415a: char_row_bitmap <= 16'b1111111111111110;
		15'h415b: char_row_bitmap <= 16'b1111111111111110;
		15'h415c: char_row_bitmap <= 16'b1111111111111110;
		15'h415d: char_row_bitmap <= 16'b1111111111111111;
		15'h415e: char_row_bitmap <= 16'b1111111111111111;
		15'h415f: char_row_bitmap <= 16'b1111111111111111;
		15'h4160: char_row_bitmap <= 16'b1111111111111111;
		15'h4161: char_row_bitmap <= 16'b1111111111111111;
		15'h4162: char_row_bitmap <= 16'b1111111111111111;
		15'h4163: char_row_bitmap <= 16'b1111111111111111;
		15'h4164: char_row_bitmap <= 16'b1111111111111111;
		15'h4165: char_row_bitmap <= 16'b1111111111111111;
		15'h4166: char_row_bitmap <= 16'b1111111111111111;
		15'h4167: char_row_bitmap <= 16'b1111111111111111;
		15'h4168: char_row_bitmap <= 16'b1111111111111111;
		15'h4169: char_row_bitmap <= 16'b1111111111111111;
		15'h416a: char_row_bitmap <= 16'b1111111111111111;
		15'h416b: char_row_bitmap <= 16'b1111111111111110;
		15'h416c: char_row_bitmap <= 16'b1111111111111110;
		15'h416d: char_row_bitmap <= 16'b1111111111111110;
		15'h416e: char_row_bitmap <= 16'b1111111111111110;
		15'h416f: char_row_bitmap <= 16'b1111111111111100;
		15'h4170: char_row_bitmap <= 16'b1111111111111100;
		15'h4171: char_row_bitmap <= 16'b1111111111111100;
		15'h4172: char_row_bitmap <= 16'b1111111111111000;
		15'h4173: char_row_bitmap <= 16'b1111111111110000;
		15'h4174: char_row_bitmap <= 16'b1111111111100000;
		15'h4175: char_row_bitmap <= 16'b1111111111000000;
		15'h4176: char_row_bitmap <= 16'b1111111100000000;
		15'h4177: char_row_bitmap <= 16'b1111000000000000;
		15'h4178: char_row_bitmap <= 16'b1111111111111111;
		15'h4179: char_row_bitmap <= 16'b1111111111111111;
		15'h417a: char_row_bitmap <= 16'b1111111111111111;
		15'h417b: char_row_bitmap <= 16'b1111111111111111;
		15'h417c: char_row_bitmap <= 16'b1111111111111111;
		15'h417d: char_row_bitmap <= 16'b1111111111111111;
		15'h417e: char_row_bitmap <= 16'b1111111111111111;
		15'h417f: char_row_bitmap <= 16'b0111111111111111;
		15'h4180: char_row_bitmap <= 16'b0111111111111111;
		15'h4181: char_row_bitmap <= 16'b0111111111111111;
		15'h4182: char_row_bitmap <= 16'b0111111111111111;
		15'h4183: char_row_bitmap <= 16'b0011111111111111;
		15'h4184: char_row_bitmap <= 16'b0011111111111111;
		15'h4185: char_row_bitmap <= 16'b0011111111111111;
		15'h4186: char_row_bitmap <= 16'b0001111111111111;
		15'h4187: char_row_bitmap <= 16'b0000111111111111;
		15'h4188: char_row_bitmap <= 16'b0000011111111111;
		15'h4189: char_row_bitmap <= 16'b0000001111111111;
		15'h418a: char_row_bitmap <= 16'b0000000011111111;
		15'h418b: char_row_bitmap <= 16'b0000000000001111;
		15'h418c: char_row_bitmap <= 16'b0000000000001111;
		15'h418d: char_row_bitmap <= 16'b0000000011111111;
		15'h418e: char_row_bitmap <= 16'b0000001111111111;
		15'h418f: char_row_bitmap <= 16'b0000011111111111;
		15'h4190: char_row_bitmap <= 16'b0000111111111111;
		15'h4191: char_row_bitmap <= 16'b0001111111111111;
		15'h4192: char_row_bitmap <= 16'b0011111111111111;
		15'h4193: char_row_bitmap <= 16'b0011111111111111;
		15'h4194: char_row_bitmap <= 16'b0011111111111111;
		15'h4195: char_row_bitmap <= 16'b0111111111111111;
		15'h4196: char_row_bitmap <= 16'b0111111111111111;
		15'h4197: char_row_bitmap <= 16'b0111111111111111;
		15'h4198: char_row_bitmap <= 16'b0111111111111111;
		15'h4199: char_row_bitmap <= 16'b1111111111111111;
		15'h419a: char_row_bitmap <= 16'b1111111111111111;
		15'h419b: char_row_bitmap <= 16'b1111111111111111;
		15'h419c: char_row_bitmap <= 16'b1111111111111111;
		15'h419d: char_row_bitmap <= 16'b1111111111111111;
		15'h419e: char_row_bitmap <= 16'b1111111111111111;
		15'h419f: char_row_bitmap <= 16'b1111111111111111;
		15'h41a0: char_row_bitmap <= 16'b0000000000000000;
		15'h41a1: char_row_bitmap <= 16'b0000000000000000;
		15'h41a2: char_row_bitmap <= 16'b0000001111000000;
		15'h41a3: char_row_bitmap <= 16'b0000111111110000;
		15'h41a4: char_row_bitmap <= 16'b0001111111111000;
		15'h41a5: char_row_bitmap <= 16'b0001111111111000;
		15'h41a6: char_row_bitmap <= 16'b0011111111111100;
		15'h41a7: char_row_bitmap <= 16'b0011111111111100;
		15'h41a8: char_row_bitmap <= 16'b0111111111111110;
		15'h41a9: char_row_bitmap <= 16'b0111111111111110;
		15'h41aa: char_row_bitmap <= 16'b0111111111111110;
		15'h41ab: char_row_bitmap <= 16'b0111111111111110;
		15'h41ac: char_row_bitmap <= 16'b0111111111111100;
		15'h41ad: char_row_bitmap <= 16'b1111111111111100;
		15'h41ae: char_row_bitmap <= 16'b1111111111111000;
		15'h41af: char_row_bitmap <= 16'b1111111111111000;
		15'h41b0: char_row_bitmap <= 16'b1111111111110000;
		15'h41b1: char_row_bitmap <= 16'b1111111111000000;
		15'h41b2: char_row_bitmap <= 16'b1111111100000000;
		15'h41b3: char_row_bitmap <= 16'b1111000000000000;
		15'h41b4: char_row_bitmap <= 16'b1111000000000000;
		15'h41b5: char_row_bitmap <= 16'b1111111100000000;
		15'h41b6: char_row_bitmap <= 16'b1111111111000000;
		15'h41b7: char_row_bitmap <= 16'b1111111111110000;
		15'h41b8: char_row_bitmap <= 16'b1111111111111000;
		15'h41b9: char_row_bitmap <= 16'b1111111111111000;
		15'h41ba: char_row_bitmap <= 16'b1111111111111100;
		15'h41bb: char_row_bitmap <= 16'b0111111111111100;
		15'h41bc: char_row_bitmap <= 16'b0111111111111110;
		15'h41bd: char_row_bitmap <= 16'b0111111111111110;
		15'h41be: char_row_bitmap <= 16'b0111111111111110;
		15'h41bf: char_row_bitmap <= 16'b0111111111111110;
		15'h41c0: char_row_bitmap <= 16'b0011111111111100;
		15'h41c1: char_row_bitmap <= 16'b0011111111111100;
		15'h41c2: char_row_bitmap <= 16'b0001111111111000;
		15'h41c3: char_row_bitmap <= 16'b0001111111111000;
		15'h41c4: char_row_bitmap <= 16'b0000111111110000;
		15'h41c5: char_row_bitmap <= 16'b0000001111000000;
		15'h41c6: char_row_bitmap <= 16'b0000000000000000;
		15'h41c7: char_row_bitmap <= 16'b0000000000000000;
		15'h41c8: char_row_bitmap <= 16'b0000000000001111;
		15'h41c9: char_row_bitmap <= 16'b0000000011111111;
		15'h41ca: char_row_bitmap <= 16'b0000001111111111;
		15'h41cb: char_row_bitmap <= 16'b0000111111111111;
		15'h41cc: char_row_bitmap <= 16'b0001111111111111;
		15'h41cd: char_row_bitmap <= 16'b0001111111111111;
		15'h41ce: char_row_bitmap <= 16'b0011111111111111;
		15'h41cf: char_row_bitmap <= 16'b0011111111111110;
		15'h41d0: char_row_bitmap <= 16'b0111111111111110;
		15'h41d1: char_row_bitmap <= 16'b0111111111111110;
		15'h41d2: char_row_bitmap <= 16'b0111111111111110;
		15'h41d3: char_row_bitmap <= 16'b0111111111111110;
		15'h41d4: char_row_bitmap <= 16'b0011111111111100;
		15'h41d5: char_row_bitmap <= 16'b0011111111111100;
		15'h41d6: char_row_bitmap <= 16'b0001111111111000;
		15'h41d7: char_row_bitmap <= 16'b0001111111111000;
		15'h41d8: char_row_bitmap <= 16'b0000111111110000;
		15'h41d9: char_row_bitmap <= 16'b0000001111000000;
		15'h41da: char_row_bitmap <= 16'b0000000000000000;
		15'h41db: char_row_bitmap <= 16'b0000000000000000;
		15'h41dc: char_row_bitmap <= 16'b0000000000000000;
		15'h41dd: char_row_bitmap <= 16'b0000000000000000;
		15'h41de: char_row_bitmap <= 16'b0000001111000000;
		15'h41df: char_row_bitmap <= 16'b0000111111110000;
		15'h41e0: char_row_bitmap <= 16'b0001111111111000;
		15'h41e1: char_row_bitmap <= 16'b0001111111111000;
		15'h41e2: char_row_bitmap <= 16'b0011111111111100;
		15'h41e3: char_row_bitmap <= 16'b0011111111111100;
		15'h41e4: char_row_bitmap <= 16'b0111111111111110;
		15'h41e5: char_row_bitmap <= 16'b0111111111111110;
		15'h41e6: char_row_bitmap <= 16'b0111111111111110;
		15'h41e7: char_row_bitmap <= 16'b0111111111111110;
		15'h41e8: char_row_bitmap <= 16'b0011111111111110;
		15'h41e9: char_row_bitmap <= 16'b0011111111111111;
		15'h41ea: char_row_bitmap <= 16'b0001111111111111;
		15'h41eb: char_row_bitmap <= 16'b0001111111111111;
		15'h41ec: char_row_bitmap <= 16'b0000111111111111;
		15'h41ed: char_row_bitmap <= 16'b0000001111111111;
		15'h41ee: char_row_bitmap <= 16'b0000000011111111;
		15'h41ef: char_row_bitmap <= 16'b0000000000001111;
		15'h41f0: char_row_bitmap <= 16'b1100000000000011;
		15'h41f1: char_row_bitmap <= 16'b1110000000000111;
		15'h41f2: char_row_bitmap <= 16'b1111000000001111;
		15'h41f3: char_row_bitmap <= 16'b1111100000011111;
		15'h41f4: char_row_bitmap <= 16'b1111100000011111;
		15'h41f5: char_row_bitmap <= 16'b1111110000111111;
		15'h41f6: char_row_bitmap <= 16'b1111110000111111;
		15'h41f7: char_row_bitmap <= 16'b1111111001111111;
		15'h41f8: char_row_bitmap <= 16'b1111111001111111;
		15'h41f9: char_row_bitmap <= 16'b1111111001111111;
		15'h41fa: char_row_bitmap <= 16'b1111111111111111;
		15'h41fb: char_row_bitmap <= 16'b1111111111111111;
		15'h41fc: char_row_bitmap <= 16'b1111111111111111;
		15'h41fd: char_row_bitmap <= 16'b1111111111111111;
		15'h41fe: char_row_bitmap <= 16'b1111111111111111;
		15'h41ff: char_row_bitmap <= 16'b1111111111111111;
		15'h4200: char_row_bitmap <= 16'b1111111111111111;
		15'h4201: char_row_bitmap <= 16'b1111111111111111;
		15'h4202: char_row_bitmap <= 16'b1111111111111111;
		15'h4203: char_row_bitmap <= 16'b1111111111111111;
		15'h4204: char_row_bitmap <= 16'b1111111111111111;
		15'h4205: char_row_bitmap <= 16'b1111111111111111;
		15'h4206: char_row_bitmap <= 16'b1111111111111110;
		15'h4207: char_row_bitmap <= 16'b1111111111111110;
		15'h4208: char_row_bitmap <= 16'b1111111111111100;
		15'h4209: char_row_bitmap <= 16'b1111111111111000;
		15'h420a: char_row_bitmap <= 16'b1111111111110000;
		15'h420b: char_row_bitmap <= 16'b1111111111000000;
		15'h420c: char_row_bitmap <= 16'b1111111100000000;
		15'h420d: char_row_bitmap <= 16'b1111110000000000;
		15'h420e: char_row_bitmap <= 16'b1111110000000000;
		15'h420f: char_row_bitmap <= 16'b1111111100000000;
		15'h4210: char_row_bitmap <= 16'b1111111111000000;
		15'h4211: char_row_bitmap <= 16'b1111111111110000;
		15'h4212: char_row_bitmap <= 16'b1111111111111000;
		15'h4213: char_row_bitmap <= 16'b1111111111111100;
		15'h4214: char_row_bitmap <= 16'b1111111111111110;
		15'h4215: char_row_bitmap <= 16'b1111111111111110;
		15'h4216: char_row_bitmap <= 16'b1111111111111111;
		15'h4217: char_row_bitmap <= 16'b1111111111111111;
		15'h4218: char_row_bitmap <= 16'b1111111111111111;
		15'h4219: char_row_bitmap <= 16'b1111111111111111;
		15'h421a: char_row_bitmap <= 16'b1111111111111111;
		15'h421b: char_row_bitmap <= 16'b1111111111111111;
		15'h421c: char_row_bitmap <= 16'b1111111111111111;
		15'h421d: char_row_bitmap <= 16'b1111111111111111;
		15'h421e: char_row_bitmap <= 16'b1111111111111111;
		15'h421f: char_row_bitmap <= 16'b1111111111111111;
		15'h4220: char_row_bitmap <= 16'b1111111111111111;
		15'h4221: char_row_bitmap <= 16'b1111111111111111;
		15'h4222: char_row_bitmap <= 16'b1111111001111111;
		15'h4223: char_row_bitmap <= 16'b1111111001111111;
		15'h4224: char_row_bitmap <= 16'b1111111001111111;
		15'h4225: char_row_bitmap <= 16'b1111110000111111;
		15'h4226: char_row_bitmap <= 16'b1111110000111111;
		15'h4227: char_row_bitmap <= 16'b1111100000011111;
		15'h4228: char_row_bitmap <= 16'b1111100000011111;
		15'h4229: char_row_bitmap <= 16'b1111000000001111;
		15'h422a: char_row_bitmap <= 16'b1110000000000111;
		15'h422b: char_row_bitmap <= 16'b1100000000000011;
		15'h422c: char_row_bitmap <= 16'b1111111111111111;
		15'h422d: char_row_bitmap <= 16'b1111111111111111;
		15'h422e: char_row_bitmap <= 16'b0111111111111111;
		15'h422f: char_row_bitmap <= 16'b0111111111111111;
		15'h4230: char_row_bitmap <= 16'b0011111111111111;
		15'h4231: char_row_bitmap <= 16'b0001111111111111;
		15'h4232: char_row_bitmap <= 16'b0000111111111111;
		15'h4233: char_row_bitmap <= 16'b0000001111111111;
		15'h4234: char_row_bitmap <= 16'b0000000011111111;
		15'h4235: char_row_bitmap <= 16'b0000000000111111;
		15'h4236: char_row_bitmap <= 16'b0000000000111111;
		15'h4237: char_row_bitmap <= 16'b0000000011111111;
		15'h4238: char_row_bitmap <= 16'b0000001111111111;
		15'h4239: char_row_bitmap <= 16'b0000111111111111;
		15'h423a: char_row_bitmap <= 16'b0001111111111111;
		15'h423b: char_row_bitmap <= 16'b0011111111111111;
		15'h423c: char_row_bitmap <= 16'b0111111111111111;
		15'h423d: char_row_bitmap <= 16'b0111111111111111;
		15'h423e: char_row_bitmap <= 16'b1111111111111111;
		15'h423f: char_row_bitmap <= 16'b1111111111111111;
		15'h4240: char_row_bitmap <= 16'b0000000000000000;
		15'h4241: char_row_bitmap <= 16'b0000000000000000;
		15'h4242: char_row_bitmap <= 16'b0000000000000000;
		15'h4243: char_row_bitmap <= 16'b0000000000000000;
		15'h4244: char_row_bitmap <= 16'b0000000000000000;
		15'h4245: char_row_bitmap <= 16'b0000000000000000;
		15'h4246: char_row_bitmap <= 16'b0000000000000000;
		15'h4247: char_row_bitmap <= 16'b0000000000000000;
		15'h4248: char_row_bitmap <= 16'b0000000000000000;
		15'h4249: char_row_bitmap <= 16'b0000000000000000;
		15'h424a: char_row_bitmap <= 16'b0000000000000000;
		15'h424b: char_row_bitmap <= 16'b0000000000000000;
		15'h424c: char_row_bitmap <= 16'b0000000000000000;
		15'h424d: char_row_bitmap <= 16'b0000000000000000;
		15'h424e: char_row_bitmap <= 16'b0000000000000000;
		15'h424f: char_row_bitmap <= 16'b0000000000000000;
		15'h4250: char_row_bitmap <= 16'b0000000000000000;
		15'h4251: char_row_bitmap <= 16'b0000000000000000;
		15'h4252: char_row_bitmap <= 16'b0000000000000000;
		15'h4253: char_row_bitmap <= 16'b0000000000000000;
		15'h4254: char_row_bitmap <= 16'b0000000000111111;
		15'h4255: char_row_bitmap <= 16'b0000000000001111;
		15'h4256: char_row_bitmap <= 16'b0000000000000011;
		15'h4257: char_row_bitmap <= 16'b0000000000000011;
		15'h4258: char_row_bitmap <= 16'b0000000000000001;
		15'h4259: char_row_bitmap <= 16'b0000000000000001;
		15'h425a: char_row_bitmap <= 16'b0000000000000000;
		15'h425b: char_row_bitmap <= 16'b0000000000000000;
		15'h425c: char_row_bitmap <= 16'b0000000000000000;
		15'h425d: char_row_bitmap <= 16'b0000000000000000;
		15'h425e: char_row_bitmap <= 16'b0000000000000000;
		15'h425f: char_row_bitmap <= 16'b0000000000000000;
		15'h4260: char_row_bitmap <= 16'b0000000000000000;
		15'h4261: char_row_bitmap <= 16'b0000000000000000;
		15'h4262: char_row_bitmap <= 16'b0000000000000000;
		15'h4263: char_row_bitmap <= 16'b0000000000000000;
		15'h4264: char_row_bitmap <= 16'b0000000000000000;
		15'h4265: char_row_bitmap <= 16'b0000000000000000;
		15'h4266: char_row_bitmap <= 16'b0000000000000000;
		15'h4267: char_row_bitmap <= 16'b0000000000000000;
		15'h4268: char_row_bitmap <= 16'b0000000000000000;
		15'h4269: char_row_bitmap <= 16'b0000000000000000;
		15'h426a: char_row_bitmap <= 16'b0000000000000000;
		15'h426b: char_row_bitmap <= 16'b0000000000000000;
		15'h426c: char_row_bitmap <= 16'b0000000000000000;
		15'h426d: char_row_bitmap <= 16'b0000000000000000;
		15'h426e: char_row_bitmap <= 16'b0000000000000000;
		15'h426f: char_row_bitmap <= 16'b0000000000000000;
		15'h4270: char_row_bitmap <= 16'b0000000000000000;
		15'h4271: char_row_bitmap <= 16'b0000000000000000;
		15'h4272: char_row_bitmap <= 16'b0000000000000000;
		15'h4273: char_row_bitmap <= 16'b0000000000000000;
		15'h4274: char_row_bitmap <= 16'b0000000000000000;
		15'h4275: char_row_bitmap <= 16'b0000000000000000;
		15'h4276: char_row_bitmap <= 16'b0000000000000001;
		15'h4277: char_row_bitmap <= 16'b0000000000000001;
		15'h4278: char_row_bitmap <= 16'b0000000000000011;
		15'h4279: char_row_bitmap <= 16'b0000000000000011;
		15'h427a: char_row_bitmap <= 16'b0000000000001111;
		15'h427b: char_row_bitmap <= 16'b0000000000111111;
		15'h427c: char_row_bitmap <= 16'b0000000000000000;
		15'h427d: char_row_bitmap <= 16'b0000000000000000;
		15'h427e: char_row_bitmap <= 16'b0000000000000000;
		15'h427f: char_row_bitmap <= 16'b0000000000000000;
		15'h4280: char_row_bitmap <= 16'b0000000000000000;
		15'h4281: char_row_bitmap <= 16'b0000000000000000;
		15'h4282: char_row_bitmap <= 16'b0000000000000000;
		15'h4283: char_row_bitmap <= 16'b0000000000000000;
		15'h4284: char_row_bitmap <= 16'b0000000000000000;
		15'h4285: char_row_bitmap <= 16'b0000000000000000;
		15'h4286: char_row_bitmap <= 16'b0000000000000000;
		15'h4287: char_row_bitmap <= 16'b0000000000000000;
		15'h4288: char_row_bitmap <= 16'b0000000000000000;
		15'h4289: char_row_bitmap <= 16'b0000000000000000;
		15'h428a: char_row_bitmap <= 16'b1000000000000000;
		15'h428b: char_row_bitmap <= 16'b1000000000000000;
		15'h428c: char_row_bitmap <= 16'b1100000000000000;
		15'h428d: char_row_bitmap <= 16'b1100000000000000;
		15'h428e: char_row_bitmap <= 16'b1111000000000000;
		15'h428f: char_row_bitmap <= 16'b1111110000000000;
		15'h4290: char_row_bitmap <= 16'b1111110000000000;
		15'h4291: char_row_bitmap <= 16'b1111000000000000;
		15'h4292: char_row_bitmap <= 16'b1100000000000000;
		15'h4293: char_row_bitmap <= 16'b1100000000000000;
		15'h4294: char_row_bitmap <= 16'b1000000000000000;
		15'h4295: char_row_bitmap <= 16'b1000000000000000;
		15'h4296: char_row_bitmap <= 16'b0000000000000000;
		15'h4297: char_row_bitmap <= 16'b0000000000000000;
		15'h4298: char_row_bitmap <= 16'b0000000000000000;
		15'h4299: char_row_bitmap <= 16'b0000000000000000;
		15'h429a: char_row_bitmap <= 16'b0000000000000000;
		15'h429b: char_row_bitmap <= 16'b0000000000000000;
		15'h429c: char_row_bitmap <= 16'b0000000000000000;
		15'h429d: char_row_bitmap <= 16'b0000000000000000;
		15'h429e: char_row_bitmap <= 16'b0000000000000000;
		15'h429f: char_row_bitmap <= 16'b0000000000000000;
		15'h42a0: char_row_bitmap <= 16'b0000000000000000;
		15'h42a1: char_row_bitmap <= 16'b0000000000000000;
		15'h42a2: char_row_bitmap <= 16'b0000000000000000;
		15'h42a3: char_row_bitmap <= 16'b0000000000000000;
		15'h42a4: char_row_bitmap <= 16'b0000000000111111;
		15'h42a5: char_row_bitmap <= 16'b0000000000001111;
		15'h42a6: char_row_bitmap <= 16'b0000000000000011;
		15'h42a7: char_row_bitmap <= 16'b0000000000000011;
		15'h42a8: char_row_bitmap <= 16'b0000000000000001;
		15'h42a9: char_row_bitmap <= 16'b0000000000000001;
		15'h42aa: char_row_bitmap <= 16'b0000000000000000;
		15'h42ab: char_row_bitmap <= 16'b0000000000000000;
		15'h42ac: char_row_bitmap <= 16'b0000000000000000;
		15'h42ad: char_row_bitmap <= 16'b0000000000000000;
		15'h42ae: char_row_bitmap <= 16'b0000000000000000;
		15'h42af: char_row_bitmap <= 16'b0000000000000000;
		15'h42b0: char_row_bitmap <= 16'b0000000000000000;
		15'h42b1: char_row_bitmap <= 16'b0000000000000000;
		15'h42b2: char_row_bitmap <= 16'b0000000000000001;
		15'h42b3: char_row_bitmap <= 16'b0000000000000001;
		15'h42b4: char_row_bitmap <= 16'b0000000000000011;
		15'h42b5: char_row_bitmap <= 16'b0000000000000011;
		15'h42b6: char_row_bitmap <= 16'b0000000000001111;
		15'h42b7: char_row_bitmap <= 16'b0000000000111111;
		15'h42b8: char_row_bitmap <= 16'b0000000000111111;
		15'h42b9: char_row_bitmap <= 16'b0000000000001111;
		15'h42ba: char_row_bitmap <= 16'b0000000000000011;
		15'h42bb: char_row_bitmap <= 16'b0000000000000011;
		15'h42bc: char_row_bitmap <= 16'b0000000000000001;
		15'h42bd: char_row_bitmap <= 16'b0000000000000001;
		15'h42be: char_row_bitmap <= 16'b0000000000000000;
		15'h42bf: char_row_bitmap <= 16'b0000000000000000;
		15'h42c0: char_row_bitmap <= 16'b0000000000000000;
		15'h42c1: char_row_bitmap <= 16'b0000000000000000;
		15'h42c2: char_row_bitmap <= 16'b0000000000000000;
		15'h42c3: char_row_bitmap <= 16'b0000000000000000;
		15'h42c4: char_row_bitmap <= 16'b0000000000000000;
		15'h42c5: char_row_bitmap <= 16'b0000000000000000;
		15'h42c6: char_row_bitmap <= 16'b1000000000000000;
		15'h42c7: char_row_bitmap <= 16'b1000000000000000;
		15'h42c8: char_row_bitmap <= 16'b1100000000000000;
		15'h42c9: char_row_bitmap <= 16'b1100000000000000;
		15'h42ca: char_row_bitmap <= 16'b1111000000000000;
		15'h42cb: char_row_bitmap <= 16'b1111110000000000;
		15'h42cc: char_row_bitmap <= 16'b1111110000111111;
		15'h42cd: char_row_bitmap <= 16'b1111000000001111;
		15'h42ce: char_row_bitmap <= 16'b1100000000000011;
		15'h42cf: char_row_bitmap <= 16'b1100000000000011;
		15'h42d0: char_row_bitmap <= 16'b1000000000000001;
		15'h42d1: char_row_bitmap <= 16'b1000000000000001;
		15'h42d2: char_row_bitmap <= 16'b0000000000000000;
		15'h42d3: char_row_bitmap <= 16'b0000000000000000;
		15'h42d4: char_row_bitmap <= 16'b0000000000000000;
		15'h42d5: char_row_bitmap <= 16'b0000000000000000;
		15'h42d6: char_row_bitmap <= 16'b0000000000000000;
		15'h42d7: char_row_bitmap <= 16'b0000000000000000;
		15'h42d8: char_row_bitmap <= 16'b0000000000000000;
		15'h42d9: char_row_bitmap <= 16'b0000000000000000;
		15'h42da: char_row_bitmap <= 16'b0000000000000000;
		15'h42db: char_row_bitmap <= 16'b0000000000000000;
		15'h42dc: char_row_bitmap <= 16'b0000000000000000;
		15'h42dd: char_row_bitmap <= 16'b0000000000000000;
		15'h42de: char_row_bitmap <= 16'b0000000000000000;
		15'h42df: char_row_bitmap <= 16'b0000000000000000;
		15'h42e0: char_row_bitmap <= 16'b0000000000000000;
		15'h42e1: char_row_bitmap <= 16'b0000000000000000;
		15'h42e2: char_row_bitmap <= 16'b0000000000000000;
		15'h42e3: char_row_bitmap <= 16'b0000000000000000;
		15'h42e4: char_row_bitmap <= 16'b0000000000000000;
		15'h42e5: char_row_bitmap <= 16'b0000000000000000;
		15'h42e6: char_row_bitmap <= 16'b0000000000000000;
		15'h42e7: char_row_bitmap <= 16'b0000000000000000;
		15'h42e8: char_row_bitmap <= 16'b0000000000000000;
		15'h42e9: char_row_bitmap <= 16'b0000000000000000;
		15'h42ea: char_row_bitmap <= 16'b0000000000000000;
		15'h42eb: char_row_bitmap <= 16'b0000000000000000;
		15'h42ec: char_row_bitmap <= 16'b0000000000000000;
		15'h42ed: char_row_bitmap <= 16'b0000000000000000;
		15'h42ee: char_row_bitmap <= 16'b1000000000000001;
		15'h42ef: char_row_bitmap <= 16'b1000000000000001;
		15'h42f0: char_row_bitmap <= 16'b1100000000000011;
		15'h42f1: char_row_bitmap <= 16'b1100000000000011;
		15'h42f2: char_row_bitmap <= 16'b1111000000001111;
		15'h42f3: char_row_bitmap <= 16'b1111110000111111;
		15'h42f4: char_row_bitmap <= 16'b1111110000000000;
		15'h42f5: char_row_bitmap <= 16'b1111000000000000;
		15'h42f6: char_row_bitmap <= 16'b1100000000000000;
		15'h42f7: char_row_bitmap <= 16'b1100000000000000;
		15'h42f8: char_row_bitmap <= 16'b1000000000000000;
		15'h42f9: char_row_bitmap <= 16'b1000000000000000;
		15'h42fa: char_row_bitmap <= 16'b0000000000000000;
		15'h42fb: char_row_bitmap <= 16'b0000000000000000;
		15'h42fc: char_row_bitmap <= 16'b0000000000000000;
		15'h42fd: char_row_bitmap <= 16'b0000000000000000;
		15'h42fe: char_row_bitmap <= 16'b0000000000000000;
		15'h42ff: char_row_bitmap <= 16'b0000000000000000;
		15'h4300: char_row_bitmap <= 16'b0000000000000000;
		15'h4301: char_row_bitmap <= 16'b0000000000000000;
		15'h4302: char_row_bitmap <= 16'b0000000000000001;
		15'h4303: char_row_bitmap <= 16'b0000000000000001;
		15'h4304: char_row_bitmap <= 16'b0000000000000011;
		15'h4305: char_row_bitmap <= 16'b0000000000000011;
		15'h4306: char_row_bitmap <= 16'b0000000000001111;
		15'h4307: char_row_bitmap <= 16'b0000000000111111;
		15'h4308: char_row_bitmap <= 16'b1111000000000000;
		15'h4309: char_row_bitmap <= 16'b1111000000000000;
		15'h430a: char_row_bitmap <= 16'b1100000000000000;
		15'h430b: char_row_bitmap <= 16'b1100000000000000;
		15'h430c: char_row_bitmap <= 16'b1000000000000000;
		15'h430d: char_row_bitmap <= 16'b1000000000000000;
		15'h430e: char_row_bitmap <= 16'b0000000000000000;
		15'h430f: char_row_bitmap <= 16'b0000000000000000;
		15'h4310: char_row_bitmap <= 16'b0000000000000000;
		15'h4311: char_row_bitmap <= 16'b0000000000000000;
		15'h4312: char_row_bitmap <= 16'b0000000000000000;
		15'h4313: char_row_bitmap <= 16'b0000000000000000;
		15'h4314: char_row_bitmap <= 16'b0000000000000000;
		15'h4315: char_row_bitmap <= 16'b0000000000000000;
		15'h4316: char_row_bitmap <= 16'b1000000000000000;
		15'h4317: char_row_bitmap <= 16'b1000000000000000;
		15'h4318: char_row_bitmap <= 16'b1100000000000000;
		15'h4319: char_row_bitmap <= 16'b1100000000000000;
		15'h431a: char_row_bitmap <= 16'b1111000000000000;
		15'h431b: char_row_bitmap <= 16'b1111110000000000;
		15'h431c: char_row_bitmap <= 16'b0000000000111111;
		15'h431d: char_row_bitmap <= 16'b0000000000001111;
		15'h431e: char_row_bitmap <= 16'b0000000000000011;
		15'h431f: char_row_bitmap <= 16'b0000000000000011;
		15'h4320: char_row_bitmap <= 16'b0000000000000001;
		15'h4321: char_row_bitmap <= 16'b0000000000000001;
		15'h4322: char_row_bitmap <= 16'b0000000000000000;
		15'h4323: char_row_bitmap <= 16'b0000000000000000;
		15'h4324: char_row_bitmap <= 16'b0000000000000000;
		15'h4325: char_row_bitmap <= 16'b0000000000000000;
		15'h4326: char_row_bitmap <= 16'b0000000000000000;
		15'h4327: char_row_bitmap <= 16'b0000000000000000;
		15'h4328: char_row_bitmap <= 16'b0000000000000000;
		15'h4329: char_row_bitmap <= 16'b0000000000000000;
		15'h432a: char_row_bitmap <= 16'b1000000000000001;
		15'h432b: char_row_bitmap <= 16'b1000000000000001;
		15'h432c: char_row_bitmap <= 16'b1100000000000011;
		15'h432d: char_row_bitmap <= 16'b1100000000000011;
		15'h432e: char_row_bitmap <= 16'b1111000000001111;
		15'h432f: char_row_bitmap <= 16'b1111110000111111;
		15'h4330: char_row_bitmap <= 16'b1111110000000000;
		15'h4331: char_row_bitmap <= 16'b1111000000000000;
		15'h4332: char_row_bitmap <= 16'b1100000000000000;
		15'h4333: char_row_bitmap <= 16'b1100000000000000;
		15'h4334: char_row_bitmap <= 16'b1000000000000000;
		15'h4335: char_row_bitmap <= 16'b1000000000000000;
		15'h4336: char_row_bitmap <= 16'b0000000000000000;
		15'h4337: char_row_bitmap <= 16'b0000000000000000;
		15'h4338: char_row_bitmap <= 16'b0000000000000000;
		15'h4339: char_row_bitmap <= 16'b0000000000000000;
		15'h433a: char_row_bitmap <= 16'b0000000000000000;
		15'h433b: char_row_bitmap <= 16'b0000000000000000;
		15'h433c: char_row_bitmap <= 16'b0000000000000000;
		15'h433d: char_row_bitmap <= 16'b0000000000000000;
		15'h433e: char_row_bitmap <= 16'b1000000000000001;
		15'h433f: char_row_bitmap <= 16'b1000000000000001;
		15'h4340: char_row_bitmap <= 16'b1100000000000011;
		15'h4341: char_row_bitmap <= 16'b1100000000000011;
		15'h4342: char_row_bitmap <= 16'b1111000000001111;
		15'h4343: char_row_bitmap <= 16'b1111110000111111;
		15'h4344: char_row_bitmap <= 16'b1111110000111111;
		15'h4345: char_row_bitmap <= 16'b1111000000001111;
		15'h4346: char_row_bitmap <= 16'b1100000000000011;
		15'h4347: char_row_bitmap <= 16'b1100000000000011;
		15'h4348: char_row_bitmap <= 16'b1000000000000001;
		15'h4349: char_row_bitmap <= 16'b1000000000000001;
		15'h434a: char_row_bitmap <= 16'b0000000000000000;
		15'h434b: char_row_bitmap <= 16'b0000000000000000;
		15'h434c: char_row_bitmap <= 16'b0000000000000000;
		15'h434d: char_row_bitmap <= 16'b0000000000000000;
		15'h434e: char_row_bitmap <= 16'b0000000000000000;
		15'h434f: char_row_bitmap <= 16'b0000000000000000;
		15'h4350: char_row_bitmap <= 16'b0000000000000000;
		15'h4351: char_row_bitmap <= 16'b0000000000000000;
		15'h4352: char_row_bitmap <= 16'b1000000000000000;
		15'h4353: char_row_bitmap <= 16'b1000000000000000;
		15'h4354: char_row_bitmap <= 16'b1100000000000000;
		15'h4355: char_row_bitmap <= 16'b1100000000000000;
		15'h4356: char_row_bitmap <= 16'b1111000000000000;
		15'h4357: char_row_bitmap <= 16'b1111110000000000;
		15'h4358: char_row_bitmap <= 16'b1111110000111111;
		15'h4359: char_row_bitmap <= 16'b1111000000001111;
		15'h435a: char_row_bitmap <= 16'b1100000000000011;
		15'h435b: char_row_bitmap <= 16'b1100000000000011;
		15'h435c: char_row_bitmap <= 16'b1000000000000001;
		15'h435d: char_row_bitmap <= 16'b1000000000000001;
		15'h435e: char_row_bitmap <= 16'b0000000000000000;
		15'h435f: char_row_bitmap <= 16'b0000000000000000;
		15'h4360: char_row_bitmap <= 16'b0000000000000000;
		15'h4361: char_row_bitmap <= 16'b0000000000000000;
		15'h4362: char_row_bitmap <= 16'b0000000000000000;
		15'h4363: char_row_bitmap <= 16'b0000000000000000;
		15'h4364: char_row_bitmap <= 16'b0000000000000000;
		15'h4365: char_row_bitmap <= 16'b0000000000000000;
		15'h4366: char_row_bitmap <= 16'b0000000000000001;
		15'h4367: char_row_bitmap <= 16'b0000000000000001;
		15'h4368: char_row_bitmap <= 16'b0000000000000011;
		15'h4369: char_row_bitmap <= 16'b0000000000000011;
		15'h436a: char_row_bitmap <= 16'b0000000000001111;
		15'h436b: char_row_bitmap <= 16'b0000000000111111;
		15'h436c: char_row_bitmap <= 16'b1111110000111111;
		15'h436d: char_row_bitmap <= 16'b1111000000001111;
		15'h436e: char_row_bitmap <= 16'b1100000000000011;
		15'h436f: char_row_bitmap <= 16'b1100000000000011;
		15'h4370: char_row_bitmap <= 16'b1000000000000001;
		15'h4371: char_row_bitmap <= 16'b1000000000000001;
		15'h4372: char_row_bitmap <= 16'b0000000000000000;
		15'h4373: char_row_bitmap <= 16'b0000000000000000;
		15'h4374: char_row_bitmap <= 16'b0000000000000000;
		15'h4375: char_row_bitmap <= 16'b0000000000000000;
		15'h4376: char_row_bitmap <= 16'b0000000000000000;
		15'h4377: char_row_bitmap <= 16'b0000000000000000;
		15'h4378: char_row_bitmap <= 16'b0000000000000000;
		15'h4379: char_row_bitmap <= 16'b0000000000000000;
		15'h437a: char_row_bitmap <= 16'b1000000000000001;
		15'h437b: char_row_bitmap <= 16'b1000000000000001;
		15'h437c: char_row_bitmap <= 16'b1100000000000011;
		15'h437d: char_row_bitmap <= 16'b1100000000000011;
		15'h437e: char_row_bitmap <= 16'b1111000000001111;
		15'h437f: char_row_bitmap <= 16'b1111110000111111;
		15'h4380: char_row_bitmap <= 16'b0000000000000000;
		15'h4381: char_row_bitmap <= 16'b0000000000000000;
		15'h4382: char_row_bitmap <= 16'b0000000000000000;
		15'h4383: char_row_bitmap <= 16'b0000000000000000;
		15'h4384: char_row_bitmap <= 16'b0011111111111111;
		15'h4385: char_row_bitmap <= 16'b0011111111111111;
		15'h4386: char_row_bitmap <= 16'b0011000000000000;
		15'h4387: char_row_bitmap <= 16'b0011000000000000;
		15'h4388: char_row_bitmap <= 16'b0011000000000000;
		15'h4389: char_row_bitmap <= 16'b0011000000000000;
		15'h438a: char_row_bitmap <= 16'b0011000000000000;
		15'h438b: char_row_bitmap <= 16'b0011000000000000;
		15'h438c: char_row_bitmap <= 16'b0011000000000000;
		15'h438d: char_row_bitmap <= 16'b0011000000000000;
		15'h438e: char_row_bitmap <= 16'b0011111111111111;
		15'h438f: char_row_bitmap <= 16'b0011111111111111;
		15'h4390: char_row_bitmap <= 16'b0000000000000000;
		15'h4391: char_row_bitmap <= 16'b0000000000000000;
		15'h4392: char_row_bitmap <= 16'b0000000000000000;
		15'h4393: char_row_bitmap <= 16'b0000000000000000;
		15'h4394: char_row_bitmap <= 16'b0000000000000000;
		15'h4395: char_row_bitmap <= 16'b0000000000000000;
		15'h4396: char_row_bitmap <= 16'b0000000000000000;
		15'h4397: char_row_bitmap <= 16'b0000000000000000;
		15'h4398: char_row_bitmap <= 16'b0011111111111111;
		15'h4399: char_row_bitmap <= 16'b0011111111111111;
		15'h439a: char_row_bitmap <= 16'b0011110000000000;
		15'h439b: char_row_bitmap <= 16'b0011110000000000;
		15'h439c: char_row_bitmap <= 16'b0011110000000000;
		15'h439d: char_row_bitmap <= 16'b0011110000000000;
		15'h439e: char_row_bitmap <= 16'b0011110000000000;
		15'h439f: char_row_bitmap <= 16'b0011110000000000;
		15'h43a0: char_row_bitmap <= 16'b0011110000000000;
		15'h43a1: char_row_bitmap <= 16'b0011110000000000;
		15'h43a2: char_row_bitmap <= 16'b0011111111111111;
		15'h43a3: char_row_bitmap <= 16'b0011111111111111;
		15'h43a4: char_row_bitmap <= 16'b0000000000000000;
		15'h43a5: char_row_bitmap <= 16'b0000000000000000;
		15'h43a6: char_row_bitmap <= 16'b0000000000000000;
		15'h43a7: char_row_bitmap <= 16'b0000000000000000;
		15'h43a8: char_row_bitmap <= 16'b0000000000000000;
		15'h43a9: char_row_bitmap <= 16'b0000000000000000;
		15'h43aa: char_row_bitmap <= 16'b0000000000000000;
		15'h43ab: char_row_bitmap <= 16'b0000000000000000;
		15'h43ac: char_row_bitmap <= 16'b0011111111111111;
		15'h43ad: char_row_bitmap <= 16'b0011111111111111;
		15'h43ae: char_row_bitmap <= 16'b0011111100000000;
		15'h43af: char_row_bitmap <= 16'b0011111100000000;
		15'h43b0: char_row_bitmap <= 16'b0011111100000000;
		15'h43b1: char_row_bitmap <= 16'b0011111100000000;
		15'h43b2: char_row_bitmap <= 16'b0011111100000000;
		15'h43b3: char_row_bitmap <= 16'b0011111100000000;
		15'h43b4: char_row_bitmap <= 16'b0011111100000000;
		15'h43b5: char_row_bitmap <= 16'b0011111100000000;
		15'h43b6: char_row_bitmap <= 16'b0011111111111111;
		15'h43b7: char_row_bitmap <= 16'b0011111111111111;
		15'h43b8: char_row_bitmap <= 16'b0000000000000000;
		15'h43b9: char_row_bitmap <= 16'b0000000000000000;
		15'h43ba: char_row_bitmap <= 16'b0000000000000000;
		15'h43bb: char_row_bitmap <= 16'b0000000000000000;
		15'h43bc: char_row_bitmap <= 16'b0000000000000000;
		15'h43bd: char_row_bitmap <= 16'b0000000000000000;
		15'h43be: char_row_bitmap <= 16'b0000000000000000;
		15'h43bf: char_row_bitmap <= 16'b0000000000000000;
		15'h43c0: char_row_bitmap <= 16'b0011111111111111;
		15'h43c1: char_row_bitmap <= 16'b0011111111111111;
		15'h43c2: char_row_bitmap <= 16'b0011111111000000;
		15'h43c3: char_row_bitmap <= 16'b0011111111000000;
		15'h43c4: char_row_bitmap <= 16'b0011111111000000;
		15'h43c5: char_row_bitmap <= 16'b0011111111000000;
		15'h43c6: char_row_bitmap <= 16'b0011111111000000;
		15'h43c7: char_row_bitmap <= 16'b0011111111000000;
		15'h43c8: char_row_bitmap <= 16'b0011111111000000;
		15'h43c9: char_row_bitmap <= 16'b0011111111000000;
		15'h43ca: char_row_bitmap <= 16'b0011111111111111;
		15'h43cb: char_row_bitmap <= 16'b0011111111111111;
		15'h43cc: char_row_bitmap <= 16'b0000000000000000;
		15'h43cd: char_row_bitmap <= 16'b0000000000000000;
		15'h43ce: char_row_bitmap <= 16'b0000000000000000;
		15'h43cf: char_row_bitmap <= 16'b0000000000000000;
		15'h43d0: char_row_bitmap <= 16'b0000000000000000;
		15'h43d1: char_row_bitmap <= 16'b0000000000000000;
		15'h43d2: char_row_bitmap <= 16'b0000000000000000;
		15'h43d3: char_row_bitmap <= 16'b0000000000000000;
		15'h43d4: char_row_bitmap <= 16'b0011111111111111;
		15'h43d5: char_row_bitmap <= 16'b0011111111111111;
		15'h43d6: char_row_bitmap <= 16'b0011111111110000;
		15'h43d7: char_row_bitmap <= 16'b0011111111110000;
		15'h43d8: char_row_bitmap <= 16'b0011111111110000;
		15'h43d9: char_row_bitmap <= 16'b0011111111110000;
		15'h43da: char_row_bitmap <= 16'b0011111111110000;
		15'h43db: char_row_bitmap <= 16'b0011111111110000;
		15'h43dc: char_row_bitmap <= 16'b0011111111110000;
		15'h43dd: char_row_bitmap <= 16'b0011111111110000;
		15'h43de: char_row_bitmap <= 16'b0011111111111111;
		15'h43df: char_row_bitmap <= 16'b0011111111111111;
		15'h43e0: char_row_bitmap <= 16'b0000000000000000;
		15'h43e1: char_row_bitmap <= 16'b0000000000000000;
		15'h43e2: char_row_bitmap <= 16'b0000000000000000;
		15'h43e3: char_row_bitmap <= 16'b0000000000000000;
		15'h43e4: char_row_bitmap <= 16'b0000000000000000;
		15'h43e5: char_row_bitmap <= 16'b0000000000000000;
		15'h43e6: char_row_bitmap <= 16'b0000000000000000;
		15'h43e7: char_row_bitmap <= 16'b0000000000000000;
		15'h43e8: char_row_bitmap <= 16'b0011111111111111;
		15'h43e9: char_row_bitmap <= 16'b0011111111111111;
		15'h43ea: char_row_bitmap <= 16'b0011111111111100;
		15'h43eb: char_row_bitmap <= 16'b0011111111111100;
		15'h43ec: char_row_bitmap <= 16'b0011111111111100;
		15'h43ed: char_row_bitmap <= 16'b0011111111111100;
		15'h43ee: char_row_bitmap <= 16'b0011111111111100;
		15'h43ef: char_row_bitmap <= 16'b0011111111111100;
		15'h43f0: char_row_bitmap <= 16'b0011111111111100;
		15'h43f1: char_row_bitmap <= 16'b0011111111111100;
		15'h43f2: char_row_bitmap <= 16'b0011111111111111;
		15'h43f3: char_row_bitmap <= 16'b0011111111111111;
		15'h43f4: char_row_bitmap <= 16'b0000000000000000;
		15'h43f5: char_row_bitmap <= 16'b0000000000000000;
		15'h43f6: char_row_bitmap <= 16'b0000000000000000;
		15'h43f7: char_row_bitmap <= 16'b0000000000000000;
		15'h43f8: char_row_bitmap <= 16'b0000000000000000;
		15'h43f9: char_row_bitmap <= 16'b0000000000000000;
		15'h43fa: char_row_bitmap <= 16'b0000000000000000;
		15'h43fb: char_row_bitmap <= 16'b0000000000000000;
		15'h43fc: char_row_bitmap <= 16'b0011111111111111;
		15'h43fd: char_row_bitmap <= 16'b0011111111111111;
		15'h43fe: char_row_bitmap <= 16'b0011111111111111;
		15'h43ff: char_row_bitmap <= 16'b0011111111111111;
		15'h4400: char_row_bitmap <= 16'b0011111111111111;
		15'h4401: char_row_bitmap <= 16'b0011111111111111;
		15'h4402: char_row_bitmap <= 16'b0011111111111111;
		15'h4403: char_row_bitmap <= 16'b0011111111111111;
		15'h4404: char_row_bitmap <= 16'b0011111111111111;
		15'h4405: char_row_bitmap <= 16'b0011111111111111;
		15'h4406: char_row_bitmap <= 16'b0011111111111111;
		15'h4407: char_row_bitmap <= 16'b0011111111111111;
		15'h4408: char_row_bitmap <= 16'b0000000000000000;
		15'h4409: char_row_bitmap <= 16'b0000000000000000;
		15'h440a: char_row_bitmap <= 16'b0000000000000000;
		15'h440b: char_row_bitmap <= 16'b0000000000000000;
		15'h440c: char_row_bitmap <= 16'b0000000000000000;
		15'h440d: char_row_bitmap <= 16'b0000000000000000;
		15'h440e: char_row_bitmap <= 16'b0000000000000000;
		15'h440f: char_row_bitmap <= 16'b0000000000000000;
		15'h4410: char_row_bitmap <= 16'b1111111111111111;
		15'h4411: char_row_bitmap <= 16'b1111111111111111;
		15'h4412: char_row_bitmap <= 16'b0000000000000000;
		15'h4413: char_row_bitmap <= 16'b0000000000000000;
		15'h4414: char_row_bitmap <= 16'b0000000000000000;
		15'h4415: char_row_bitmap <= 16'b0000000000000000;
		15'h4416: char_row_bitmap <= 16'b0000000000000000;
		15'h4417: char_row_bitmap <= 16'b0000000000000000;
		15'h4418: char_row_bitmap <= 16'b0000000000000000;
		15'h4419: char_row_bitmap <= 16'b0000000000000000;
		15'h441a: char_row_bitmap <= 16'b1111111111111111;
		15'h441b: char_row_bitmap <= 16'b1111111111111111;
		15'h441c: char_row_bitmap <= 16'b0000000000000000;
		15'h441d: char_row_bitmap <= 16'b0000000000000000;
		15'h441e: char_row_bitmap <= 16'b0000000000000000;
		15'h441f: char_row_bitmap <= 16'b0000000000000000;
		15'h4420: char_row_bitmap <= 16'b0000000000000000;
		15'h4421: char_row_bitmap <= 16'b0000000000000000;
		15'h4422: char_row_bitmap <= 16'b0000000000000000;
		15'h4423: char_row_bitmap <= 16'b0000000000000000;
		15'h4424: char_row_bitmap <= 16'b1111111111111111;
		15'h4425: char_row_bitmap <= 16'b1111111111111111;
		15'h4426: char_row_bitmap <= 16'b1100000000000000;
		15'h4427: char_row_bitmap <= 16'b1100000000000000;
		15'h4428: char_row_bitmap <= 16'b1100000000000000;
		15'h4429: char_row_bitmap <= 16'b1100000000000000;
		15'h442a: char_row_bitmap <= 16'b1100000000000000;
		15'h442b: char_row_bitmap <= 16'b1100000000000000;
		15'h442c: char_row_bitmap <= 16'b1100000000000000;
		15'h442d: char_row_bitmap <= 16'b1100000000000000;
		15'h442e: char_row_bitmap <= 16'b1111111111111111;
		15'h442f: char_row_bitmap <= 16'b1111111111111111;
		15'h4430: char_row_bitmap <= 16'b0000000000000000;
		15'h4431: char_row_bitmap <= 16'b0000000000000000;
		15'h4432: char_row_bitmap <= 16'b0000000000000000;
		15'h4433: char_row_bitmap <= 16'b0000000000000000;
		15'h4434: char_row_bitmap <= 16'b0000000000000000;
		15'h4435: char_row_bitmap <= 16'b0000000000000000;
		15'h4436: char_row_bitmap <= 16'b0000000000000000;
		15'h4437: char_row_bitmap <= 16'b0000000000000000;
		15'h4438: char_row_bitmap <= 16'b1111111111111111;
		15'h4439: char_row_bitmap <= 16'b1111111111111111;
		15'h443a: char_row_bitmap <= 16'b1111000000000000;
		15'h443b: char_row_bitmap <= 16'b1111000000000000;
		15'h443c: char_row_bitmap <= 16'b1111000000000000;
		15'h443d: char_row_bitmap <= 16'b1111000000000000;
		15'h443e: char_row_bitmap <= 16'b1111000000000000;
		15'h443f: char_row_bitmap <= 16'b1111000000000000;
		15'h4440: char_row_bitmap <= 16'b1111000000000000;
		15'h4441: char_row_bitmap <= 16'b1111000000000000;
		15'h4442: char_row_bitmap <= 16'b1111111111111111;
		15'h4443: char_row_bitmap <= 16'b1111111111111111;
		15'h4444: char_row_bitmap <= 16'b0000000000000000;
		15'h4445: char_row_bitmap <= 16'b0000000000000000;
		15'h4446: char_row_bitmap <= 16'b0000000000000000;
		15'h4447: char_row_bitmap <= 16'b0000000000000000;
		15'h4448: char_row_bitmap <= 16'b0000000000000000;
		15'h4449: char_row_bitmap <= 16'b0000000000000000;
		15'h444a: char_row_bitmap <= 16'b0000000000000000;
		15'h444b: char_row_bitmap <= 16'b0000000000000000;
		15'h444c: char_row_bitmap <= 16'b1111111111111111;
		15'h444d: char_row_bitmap <= 16'b1111111111111111;
		15'h444e: char_row_bitmap <= 16'b1111110000000000;
		15'h444f: char_row_bitmap <= 16'b1111110000000000;
		15'h4450: char_row_bitmap <= 16'b1111110000000000;
		15'h4451: char_row_bitmap <= 16'b1111110000000000;
		15'h4452: char_row_bitmap <= 16'b1111110000000000;
		15'h4453: char_row_bitmap <= 16'b1111110000000000;
		15'h4454: char_row_bitmap <= 16'b1111110000000000;
		15'h4455: char_row_bitmap <= 16'b1111110000000000;
		15'h4456: char_row_bitmap <= 16'b1111111111111111;
		15'h4457: char_row_bitmap <= 16'b1111111111111111;
		15'h4458: char_row_bitmap <= 16'b0000000000000000;
		15'h4459: char_row_bitmap <= 16'b0000000000000000;
		15'h445a: char_row_bitmap <= 16'b0000000000000000;
		15'h445b: char_row_bitmap <= 16'b0000000000000000;
		15'h445c: char_row_bitmap <= 16'b0000000000000000;
		15'h445d: char_row_bitmap <= 16'b0000000000000000;
		15'h445e: char_row_bitmap <= 16'b0000000000000000;
		15'h445f: char_row_bitmap <= 16'b0000000000000000;
		15'h4460: char_row_bitmap <= 16'b1111111111111111;
		15'h4461: char_row_bitmap <= 16'b1111111111111111;
		15'h4462: char_row_bitmap <= 16'b1111111100000000;
		15'h4463: char_row_bitmap <= 16'b1111111100000000;
		15'h4464: char_row_bitmap <= 16'b1111111100000000;
		15'h4465: char_row_bitmap <= 16'b1111111100000000;
		15'h4466: char_row_bitmap <= 16'b1111111100000000;
		15'h4467: char_row_bitmap <= 16'b1111111100000000;
		15'h4468: char_row_bitmap <= 16'b1111111100000000;
		15'h4469: char_row_bitmap <= 16'b1111111100000000;
		15'h446a: char_row_bitmap <= 16'b1111111111111111;
		15'h446b: char_row_bitmap <= 16'b1111111111111111;
		15'h446c: char_row_bitmap <= 16'b0000000000000000;
		15'h446d: char_row_bitmap <= 16'b0000000000000000;
		15'h446e: char_row_bitmap <= 16'b0000000000000000;
		15'h446f: char_row_bitmap <= 16'b0000000000000000;
		15'h4470: char_row_bitmap <= 16'b0000000000000000;
		15'h4471: char_row_bitmap <= 16'b0000000000000000;
		15'h4472: char_row_bitmap <= 16'b0000000000000000;
		15'h4473: char_row_bitmap <= 16'b0000000000000000;
		15'h4474: char_row_bitmap <= 16'b1111111111111111;
		15'h4475: char_row_bitmap <= 16'b1111111111111111;
		15'h4476: char_row_bitmap <= 16'b1111111111000000;
		15'h4477: char_row_bitmap <= 16'b1111111111000000;
		15'h4478: char_row_bitmap <= 16'b1111111111000000;
		15'h4479: char_row_bitmap <= 16'b1111111111000000;
		15'h447a: char_row_bitmap <= 16'b1111111111000000;
		15'h447b: char_row_bitmap <= 16'b1111111111000000;
		15'h447c: char_row_bitmap <= 16'b1111111111000000;
		15'h447d: char_row_bitmap <= 16'b1111111111000000;
		15'h447e: char_row_bitmap <= 16'b1111111111111111;
		15'h447f: char_row_bitmap <= 16'b1111111111111111;
		15'h4480: char_row_bitmap <= 16'b0000000000000000;
		15'h4481: char_row_bitmap <= 16'b0000000000000000;
		15'h4482: char_row_bitmap <= 16'b0000000000000000;
		15'h4483: char_row_bitmap <= 16'b0000000000000000;
		15'h4484: char_row_bitmap <= 16'b0000000000000000;
		15'h4485: char_row_bitmap <= 16'b0000000000000000;
		15'h4486: char_row_bitmap <= 16'b0000000000000000;
		15'h4487: char_row_bitmap <= 16'b0000000000000000;
		15'h4488: char_row_bitmap <= 16'b1111111111111111;
		15'h4489: char_row_bitmap <= 16'b1111111111111111;
		15'h448a: char_row_bitmap <= 16'b1111111111110000;
		15'h448b: char_row_bitmap <= 16'b1111111111110000;
		15'h448c: char_row_bitmap <= 16'b1111111111110000;
		15'h448d: char_row_bitmap <= 16'b1111111111110000;
		15'h448e: char_row_bitmap <= 16'b1111111111110000;
		15'h448f: char_row_bitmap <= 16'b1111111111110000;
		15'h4490: char_row_bitmap <= 16'b1111111111110000;
		15'h4491: char_row_bitmap <= 16'b1111111111110000;
		15'h4492: char_row_bitmap <= 16'b1111111111111111;
		15'h4493: char_row_bitmap <= 16'b1111111111111111;
		15'h4494: char_row_bitmap <= 16'b0000000000000000;
		15'h4495: char_row_bitmap <= 16'b0000000000000000;
		15'h4496: char_row_bitmap <= 16'b0000000000000000;
		15'h4497: char_row_bitmap <= 16'b0000000000000000;
		15'h4498: char_row_bitmap <= 16'b0000000000000000;
		15'h4499: char_row_bitmap <= 16'b0000000000000000;
		15'h449a: char_row_bitmap <= 16'b0000000000000000;
		15'h449b: char_row_bitmap <= 16'b0000000000000000;
		15'h449c: char_row_bitmap <= 16'b1111111111111111;
		15'h449d: char_row_bitmap <= 16'b1111111111111111;
		15'h449e: char_row_bitmap <= 16'b1111111111111100;
		15'h449f: char_row_bitmap <= 16'b1111111111111100;
		15'h44a0: char_row_bitmap <= 16'b1111111111111100;
		15'h44a1: char_row_bitmap <= 16'b1111111111111100;
		15'h44a2: char_row_bitmap <= 16'b1111111111111100;
		15'h44a3: char_row_bitmap <= 16'b1111111111111100;
		15'h44a4: char_row_bitmap <= 16'b1111111111111100;
		15'h44a5: char_row_bitmap <= 16'b1111111111111100;
		15'h44a6: char_row_bitmap <= 16'b1111111111111111;
		15'h44a7: char_row_bitmap <= 16'b1111111111111111;
		15'h44a8: char_row_bitmap <= 16'b0000000000000000;
		15'h44a9: char_row_bitmap <= 16'b0000000000000000;
		15'h44aa: char_row_bitmap <= 16'b0000000000000000;
		15'h44ab: char_row_bitmap <= 16'b0000000000000000;
		15'h44ac: char_row_bitmap <= 16'b0000000000000000;
		15'h44ad: char_row_bitmap <= 16'b0000000000000000;
		15'h44ae: char_row_bitmap <= 16'b0000000000000000;
		15'h44af: char_row_bitmap <= 16'b0000000000000000;
		15'h44b0: char_row_bitmap <= 16'b1111111111111111;
		15'h44b1: char_row_bitmap <= 16'b1111111111111111;
		15'h44b2: char_row_bitmap <= 16'b1111111111111111;
		15'h44b3: char_row_bitmap <= 16'b1111111111111111;
		15'h44b4: char_row_bitmap <= 16'b1111111111111111;
		15'h44b5: char_row_bitmap <= 16'b1111111111111111;
		15'h44b6: char_row_bitmap <= 16'b1111111111111111;
		15'h44b7: char_row_bitmap <= 16'b1111111111111111;
		15'h44b8: char_row_bitmap <= 16'b1111111111111111;
		15'h44b9: char_row_bitmap <= 16'b1111111111111111;
		15'h44ba: char_row_bitmap <= 16'b1111111111111111;
		15'h44bb: char_row_bitmap <= 16'b1111111111111111;
		15'h44bc: char_row_bitmap <= 16'b0000000000000000;
		15'h44bd: char_row_bitmap <= 16'b0000000000000000;
		15'h44be: char_row_bitmap <= 16'b0000000000000000;
		15'h44bf: char_row_bitmap <= 16'b0000000000000000;
		15'h44c0: char_row_bitmap <= 16'b0000000000000000;
		15'h44c1: char_row_bitmap <= 16'b0000000000000000;
		15'h44c2: char_row_bitmap <= 16'b0000000000000000;
		15'h44c3: char_row_bitmap <= 16'b0000000000000000;
		15'h44c4: char_row_bitmap <= 16'b1111111111110000;
		15'h44c5: char_row_bitmap <= 16'b1111111111110000;
		15'h44c6: char_row_bitmap <= 16'b0000000000110000;
		15'h44c7: char_row_bitmap <= 16'b0000000000110000;
		15'h44c8: char_row_bitmap <= 16'b0000000000110000;
		15'h44c9: char_row_bitmap <= 16'b0000000000110000;
		15'h44ca: char_row_bitmap <= 16'b0000000000110000;
		15'h44cb: char_row_bitmap <= 16'b0000000000110000;
		15'h44cc: char_row_bitmap <= 16'b0000000000110000;
		15'h44cd: char_row_bitmap <= 16'b0000000000110000;
		15'h44ce: char_row_bitmap <= 16'b1111111111110000;
		15'h44cf: char_row_bitmap <= 16'b1111111111110000;
		15'h44d0: char_row_bitmap <= 16'b0000000000000000;
		15'h44d1: char_row_bitmap <= 16'b0000000000000000;
		15'h44d2: char_row_bitmap <= 16'b0000000000000000;
		15'h44d3: char_row_bitmap <= 16'b0000000000000000;
		15'h44d4: char_row_bitmap <= 16'b0000000000000000;
		15'h44d5: char_row_bitmap <= 16'b0000000000000000;
		15'h44d6: char_row_bitmap <= 16'b0000000000000000;
		15'h44d7: char_row_bitmap <= 16'b0000000000000000;
		15'h44d8: char_row_bitmap <= 16'b1111111111110000;
		15'h44d9: char_row_bitmap <= 16'b1111111111110000;
		15'h44da: char_row_bitmap <= 16'b1100000000110000;
		15'h44db: char_row_bitmap <= 16'b1100000000110000;
		15'h44dc: char_row_bitmap <= 16'b1100000000110000;
		15'h44dd: char_row_bitmap <= 16'b1100000000110000;
		15'h44de: char_row_bitmap <= 16'b1100000000110000;
		15'h44df: char_row_bitmap <= 16'b1100000000110000;
		15'h44e0: char_row_bitmap <= 16'b1100000000110000;
		15'h44e1: char_row_bitmap <= 16'b1100000000110000;
		15'h44e2: char_row_bitmap <= 16'b1111111111110000;
		15'h44e3: char_row_bitmap <= 16'b1111111111110000;
		15'h44e4: char_row_bitmap <= 16'b0000000000000000;
		15'h44e5: char_row_bitmap <= 16'b0000000000000000;
		15'h44e6: char_row_bitmap <= 16'b0000000000000000;
		15'h44e7: char_row_bitmap <= 16'b0000000000000000;
		15'h44e8: char_row_bitmap <= 16'b0000000000000000;
		15'h44e9: char_row_bitmap <= 16'b0000000000000000;
		15'h44ea: char_row_bitmap <= 16'b0000000000000000;
		15'h44eb: char_row_bitmap <= 16'b0000000000000000;
		15'h44ec: char_row_bitmap <= 16'b1111111111110000;
		15'h44ed: char_row_bitmap <= 16'b1111111111110000;
		15'h44ee: char_row_bitmap <= 16'b1111000000110000;
		15'h44ef: char_row_bitmap <= 16'b1111000000110000;
		15'h44f0: char_row_bitmap <= 16'b1111000000110000;
		15'h44f1: char_row_bitmap <= 16'b1111000000110000;
		15'h44f2: char_row_bitmap <= 16'b1111000000110000;
		15'h44f3: char_row_bitmap <= 16'b1111000000110000;
		15'h44f4: char_row_bitmap <= 16'b1111000000110000;
		15'h44f5: char_row_bitmap <= 16'b1111000000110000;
		15'h44f6: char_row_bitmap <= 16'b1111111111110000;
		15'h44f7: char_row_bitmap <= 16'b1111111111110000;
		15'h44f8: char_row_bitmap <= 16'b0000000000000000;
		15'h44f9: char_row_bitmap <= 16'b0000000000000000;
		15'h44fa: char_row_bitmap <= 16'b0000000000000000;
		15'h44fb: char_row_bitmap <= 16'b0000000000000000;
		15'h44fc: char_row_bitmap <= 16'b0000000000000000;
		15'h44fd: char_row_bitmap <= 16'b0000000000000000;
		15'h44fe: char_row_bitmap <= 16'b0000000000000000;
		15'h44ff: char_row_bitmap <= 16'b0000000000000000;
		15'h4500: char_row_bitmap <= 16'b1111111111110000;
		15'h4501: char_row_bitmap <= 16'b1111111111110000;
		15'h4502: char_row_bitmap <= 16'b1111110000110000;
		15'h4503: char_row_bitmap <= 16'b1111110000110000;
		15'h4504: char_row_bitmap <= 16'b1111110000110000;
		15'h4505: char_row_bitmap <= 16'b1111110000110000;
		15'h4506: char_row_bitmap <= 16'b1111110000110000;
		15'h4507: char_row_bitmap <= 16'b1111110000110000;
		15'h4508: char_row_bitmap <= 16'b1111110000110000;
		15'h4509: char_row_bitmap <= 16'b1111110000110000;
		15'h450a: char_row_bitmap <= 16'b1111111111110000;
		15'h450b: char_row_bitmap <= 16'b1111111111110000;
		15'h450c: char_row_bitmap <= 16'b0000000000000000;
		15'h450d: char_row_bitmap <= 16'b0000000000000000;
		15'h450e: char_row_bitmap <= 16'b0000000000000000;
		15'h450f: char_row_bitmap <= 16'b0000000000000000;
		15'h4510: char_row_bitmap <= 16'b0000000000000000;
		15'h4511: char_row_bitmap <= 16'b0000000000000000;
		15'h4512: char_row_bitmap <= 16'b0000000000000000;
		15'h4513: char_row_bitmap <= 16'b0000000000000000;
		15'h4514: char_row_bitmap <= 16'b1111111111110000;
		15'h4515: char_row_bitmap <= 16'b1111111111110000;
		15'h4516: char_row_bitmap <= 16'b1111111100110000;
		15'h4517: char_row_bitmap <= 16'b1111111100110000;
		15'h4518: char_row_bitmap <= 16'b1111111100110000;
		15'h4519: char_row_bitmap <= 16'b1111111100110000;
		15'h451a: char_row_bitmap <= 16'b1111111100110000;
		15'h451b: char_row_bitmap <= 16'b1111111100110000;
		15'h451c: char_row_bitmap <= 16'b1111111100110000;
		15'h451d: char_row_bitmap <= 16'b1111111100110000;
		15'h451e: char_row_bitmap <= 16'b1111111111110000;
		15'h451f: char_row_bitmap <= 16'b1111111111110000;
		15'h4520: char_row_bitmap <= 16'b0000000000000000;
		15'h4521: char_row_bitmap <= 16'b0000000000000000;
		15'h4522: char_row_bitmap <= 16'b0000000000000000;
		15'h4523: char_row_bitmap <= 16'b0000000000000000;
		15'h4524: char_row_bitmap <= 16'b0000000000000000;
		15'h4525: char_row_bitmap <= 16'b0000000000000000;
		15'h4526: char_row_bitmap <= 16'b0000000000000000;
		15'h4527: char_row_bitmap <= 16'b0000000000000000;
		15'h4528: char_row_bitmap <= 16'b1111111111110000;
		15'h4529: char_row_bitmap <= 16'b1111111111110000;
		15'h452a: char_row_bitmap <= 16'b1111111111110000;
		15'h452b: char_row_bitmap <= 16'b1111111111110000;
		15'h452c: char_row_bitmap <= 16'b1111111111110000;
		15'h452d: char_row_bitmap <= 16'b1111111111110000;
		15'h452e: char_row_bitmap <= 16'b1111111111110000;
		15'h452f: char_row_bitmap <= 16'b1111111111110000;
		15'h4530: char_row_bitmap <= 16'b1111111111110000;
		15'h4531: char_row_bitmap <= 16'b1111111111110000;
		15'h4532: char_row_bitmap <= 16'b1111111111110000;
		15'h4533: char_row_bitmap <= 16'b1111111111110000;
		15'h4534: char_row_bitmap <= 16'b0000000000000000;
		15'h4535: char_row_bitmap <= 16'b0000000000000000;
		15'h4536: char_row_bitmap <= 16'b0000000000000000;
		15'h4537: char_row_bitmap <= 16'b0000000000000000;
		15'h4538: char_row_bitmap <= 16'b0000000000000000;
		15'h4539: char_row_bitmap <= 16'b0000000000000000;
		15'h453a: char_row_bitmap <= 16'b0000000000000000;
		15'h453b: char_row_bitmap <= 16'b0000000000000000;
		15'h453c: char_row_bitmap <= 16'b0000000000000000;
		15'h453d: char_row_bitmap <= 16'b0000001111111100;
		15'h453e: char_row_bitmap <= 16'b0000010000000100;
		15'h453f: char_row_bitmap <= 16'b0000100100010100;
		15'h4540: char_row_bitmap <= 16'b0001000010100100;
		15'h4541: char_row_bitmap <= 16'b0010000001000100;
		15'h4542: char_row_bitmap <= 16'b0001000010100100;
		15'h4543: char_row_bitmap <= 16'b0000100100010100;
		15'h4544: char_row_bitmap <= 16'b0000010000000100;
		15'h4545: char_row_bitmap <= 16'b0000001111111100;
		15'h4546: char_row_bitmap <= 16'b0000000000000000;
		15'h4547: char_row_bitmap <= 16'b0000000000000000;
		15'h4548: char_row_bitmap <= 16'b0000000000000000;
		15'h4549: char_row_bitmap <= 16'b0000000000000000;
		15'h454a: char_row_bitmap <= 16'b0000000000000000;
		15'h454b: char_row_bitmap <= 16'b0000000000000000;
		15'h454c: char_row_bitmap <= 16'b0000000000000000;
		15'h454d: char_row_bitmap <= 16'b0000000000000000;
		15'h454e: char_row_bitmap <= 16'b0000000000000000;
		15'h454f: char_row_bitmap <= 16'b0000000000000000;
		15'h4550: char_row_bitmap <= 16'b0000000000000000;
		15'h4551: char_row_bitmap <= 16'b0011111111000000;
		15'h4552: char_row_bitmap <= 16'b0010000000100000;
		15'h4553: char_row_bitmap <= 16'b0010100010010000;
		15'h4554: char_row_bitmap <= 16'b0010010100001000;
		15'h4555: char_row_bitmap <= 16'b0010001000000100;
		15'h4556: char_row_bitmap <= 16'b0010010100001000;
		15'h4557: char_row_bitmap <= 16'b0010100010010000;
		15'h4558: char_row_bitmap <= 16'b0010000000100000;
		15'h4559: char_row_bitmap <= 16'b0011111111000000;
		15'h455a: char_row_bitmap <= 16'b0000000000000000;
		15'h455b: char_row_bitmap <= 16'b0000000000000000;
		15'h455c: char_row_bitmap <= 16'b0000000000000000;
		15'h455d: char_row_bitmap <= 16'b0000000000000000;
		15'h455e: char_row_bitmap <= 16'b0000000000000000;
		15'h455f: char_row_bitmap <= 16'b0000000000000000;
		15'h4560: char_row_bitmap <= 16'b0000000000000000;
		15'h4561: char_row_bitmap <= 16'b0000000000000000;
		15'h4562: char_row_bitmap <= 16'b0000000110000000;
		15'h4563: char_row_bitmap <= 16'b0000011111100000;
		15'h4564: char_row_bitmap <= 16'b0000111111110000;
		15'h4565: char_row_bitmap <= 16'b0001110000111000;
		15'h4566: char_row_bitmap <= 16'b0001100000011000;
		15'h4567: char_row_bitmap <= 16'b0001100000011000;
		15'h4568: char_row_bitmap <= 16'b0001100000011000;
		15'h4569: char_row_bitmap <= 16'b0011111111111100;
		15'h456a: char_row_bitmap <= 16'b0011111111111100;
		15'h456b: char_row_bitmap <= 16'b0011000000001100;
		15'h456c: char_row_bitmap <= 16'b0011001111001100;
		15'h456d: char_row_bitmap <= 16'b0011001111001100;
		15'h456e: char_row_bitmap <= 16'b0011000110001100;
		15'h456f: char_row_bitmap <= 16'b0011000110001100;
		15'h4570: char_row_bitmap <= 16'b0011000000001100;
		15'h4571: char_row_bitmap <= 16'b0011111111111100;
		15'h4572: char_row_bitmap <= 16'b0011111111111100;
		15'h4573: char_row_bitmap <= 16'b0000000000000000;
		15'h4574: char_row_bitmap <= 16'b0000000000000000;
		15'h4575: char_row_bitmap <= 16'b0000000000000000;
		15'h4576: char_row_bitmap <= 16'b0000000000000000;
		15'h4577: char_row_bitmap <= 16'b0000000000000000;
		15'h4578: char_row_bitmap <= 16'b0000000000000000;
		15'h4579: char_row_bitmap <= 16'b0000000000000000;
		15'h457a: char_row_bitmap <= 16'b0000000000000000;
		15'h457b: char_row_bitmap <= 16'b0000000000000000;
		15'h457c: char_row_bitmap <= 16'b0000000000000000;
		15'h457d: char_row_bitmap <= 16'b0000000000000000;
		15'h457e: char_row_bitmap <= 16'b0000000000000000;
		15'h457f: char_row_bitmap <= 16'b0000000000000000;
		15'h4580: char_row_bitmap <= 16'b0000000000000000;
		15'h4581: char_row_bitmap <= 16'b0000000000000000;
		15'h4582: char_row_bitmap <= 16'b0000000000000000;
		15'h4583: char_row_bitmap <= 16'b0000000000000000;
		15'h4584: char_row_bitmap <= 16'b0000000000000000;
		15'h4585: char_row_bitmap <= 16'b0000000000000000;
		15'h4586: char_row_bitmap <= 16'b0000000000000000;
		15'h4587: char_row_bitmap <= 16'b0000000000000000;
		15'h4588: char_row_bitmap <= 16'b0000000000000000;
		15'h4589: char_row_bitmap <= 16'b0000000000000000;
		15'h458a: char_row_bitmap <= 16'b0000000000000000;
		15'h458b: char_row_bitmap <= 16'b0000000000000000;
		15'h458c: char_row_bitmap <= 16'b0000000000000000;
		15'h458d: char_row_bitmap <= 16'b0000000000000000;
		15'h458e: char_row_bitmap <= 16'b0000000000000000;
		15'h458f: char_row_bitmap <= 16'b0000000000000000;
		15'h4590: char_row_bitmap <= 16'b0000000000000000;
		15'h4591: char_row_bitmap <= 16'b0000000000000000;
		15'h4592: char_row_bitmap <= 16'b0000000000000000;
		15'h4593: char_row_bitmap <= 16'b0000000000000000;
		15'h4594: char_row_bitmap <= 16'b0000000000000000;
		15'h4595: char_row_bitmap <= 16'b0000000000000000;
		15'h4596: char_row_bitmap <= 16'b0000000000000000;
		15'h4597: char_row_bitmap <= 16'b0000000000000000;
		15'h4598: char_row_bitmap <= 16'b0000000000000000;
		15'h4599: char_row_bitmap <= 16'b0000000000000000;
		15'h459a: char_row_bitmap <= 16'b0000000000000000;
		15'h459b: char_row_bitmap <= 16'b0000000000000000;
		15'h459c: char_row_bitmap <= 16'b0000000000000000;
		15'h459d: char_row_bitmap <= 16'b0000000000000000;
		15'h459e: char_row_bitmap <= 16'b0000000000000000;
		15'h459f: char_row_bitmap <= 16'b0000000000000000;
		15'h45a0: char_row_bitmap <= 16'b0000000000000000;
		15'h45a1: char_row_bitmap <= 16'b0000000000000000;
		15'h45a2: char_row_bitmap <= 16'b0000000000000000;
		15'h45a3: char_row_bitmap <= 16'b0000000000000000;
		15'h45a4: char_row_bitmap <= 16'b0000000000000000;
		15'h45a5: char_row_bitmap <= 16'b0000000000000000;
		15'h45a6: char_row_bitmap <= 16'b0000000000000000;
		15'h45a7: char_row_bitmap <= 16'b0000000000000000;
		15'h45a8: char_row_bitmap <= 16'b0000000000000000;
		15'h45a9: char_row_bitmap <= 16'b0000000000000000;
		15'h45aa: char_row_bitmap <= 16'b0000000000000000;
		15'h45ab: char_row_bitmap <= 16'b0000000000000000;
		15'h45ac: char_row_bitmap <= 16'b0000000000000000;
		15'h45ad: char_row_bitmap <= 16'b0000000000000000;
		15'h45ae: char_row_bitmap <= 16'b0000000000000000;
		15'h45af: char_row_bitmap <= 16'b0000000000000000;
		15'h45b0: char_row_bitmap <= 16'b0000000000000000;
		15'h45b1: char_row_bitmap <= 16'b0000000000000000;
		15'h45b2: char_row_bitmap <= 16'b0000000000000000;
		15'h45b3: char_row_bitmap <= 16'b0000000000000000;
		15'h45b4: char_row_bitmap <= 16'b0000000000000000;
		15'h45b5: char_row_bitmap <= 16'b0000000000000000;
		15'h45b6: char_row_bitmap <= 16'b0000000000000000;
		15'h45b7: char_row_bitmap <= 16'b0000000000000000;
		15'h45b8: char_row_bitmap <= 16'b0000000000000000;
		15'h45b9: char_row_bitmap <= 16'b0000000000000000;
		15'h45ba: char_row_bitmap <= 16'b0000000000000000;
		15'h45bb: char_row_bitmap <= 16'b0000000000000000;
		15'h45bc: char_row_bitmap <= 16'b0000000000000000;
		15'h45bd: char_row_bitmap <= 16'b0000000000000000;
		15'h45be: char_row_bitmap <= 16'b0000000000000000;
		15'h45bf: char_row_bitmap <= 16'b0000000000000000;
		15'h45c0: char_row_bitmap <= 16'b0000000000000000;
		15'h45c1: char_row_bitmap <= 16'b0000000000000000;
		15'h45c2: char_row_bitmap <= 16'b0000000000000000;
		15'h45c3: char_row_bitmap <= 16'b0000000000000000;
		15'h45c4: char_row_bitmap <= 16'b0000000000000000;
		15'h45c5: char_row_bitmap <= 16'b0000000000000000;
		15'h45c6: char_row_bitmap <= 16'b0000000000000000;
		15'h45c7: char_row_bitmap <= 16'b0000000000000000;
		15'h45c8: char_row_bitmap <= 16'b0000000000000000;
		15'h45c9: char_row_bitmap <= 16'b0000000000000000;
		15'h45ca: char_row_bitmap <= 16'b0000000000000000;
		15'h45cb: char_row_bitmap <= 16'b0000000000000000;
		15'h45cc: char_row_bitmap <= 16'b0000000000000000;
		15'h45cd: char_row_bitmap <= 16'b0000000000000000;
		15'h45ce: char_row_bitmap <= 16'b0000000000000000;
		15'h45cf: char_row_bitmap <= 16'b0000000000000000;
		15'h45d0: char_row_bitmap <= 16'b0000000000000000;
		15'h45d1: char_row_bitmap <= 16'b0000000000000000;
		15'h45d2: char_row_bitmap <= 16'b0000000000000000;
		15'h45d3: char_row_bitmap <= 16'b0000000000000000;
		15'h45d4: char_row_bitmap <= 16'b0000000000000000;
		15'h45d5: char_row_bitmap <= 16'b0000000000000000;
		15'h45d6: char_row_bitmap <= 16'b0000000000000000;
		15'h45d7: char_row_bitmap <= 16'b0000000000000000;
		15'h45d8: char_row_bitmap <= 16'b0000000000000000;
		15'h45d9: char_row_bitmap <= 16'b0000000000000000;
		15'h45da: char_row_bitmap <= 16'b0000000000000000;
		15'h45db: char_row_bitmap <= 16'b0000000000000000;
		15'h45dc: char_row_bitmap <= 16'b0000000000000000;
		15'h45dd: char_row_bitmap <= 16'b0000000000000000;
		15'h45de: char_row_bitmap <= 16'b0000000000000000;
		15'h45df: char_row_bitmap <= 16'b0000000000000000;
		15'h45e0: char_row_bitmap <= 16'b0000000000000000;
		15'h45e1: char_row_bitmap <= 16'b0000000000000000;
		15'h45e2: char_row_bitmap <= 16'b0000000000000000;
		15'h45e3: char_row_bitmap <= 16'b0000000000000000;
		15'h45e4: char_row_bitmap <= 16'b0000000000000000;
		15'h45e5: char_row_bitmap <= 16'b0000000000000000;
		15'h45e6: char_row_bitmap <= 16'b0000000000000000;
		15'h45e7: char_row_bitmap <= 16'b0000000000000000;
		15'h45e8: char_row_bitmap <= 16'b0000000000000000;
		15'h45e9: char_row_bitmap <= 16'b0000000000000000;
		15'h45ea: char_row_bitmap <= 16'b0000000000000000;
		15'h45eb: char_row_bitmap <= 16'b0000000000000000;
		15'h45ec: char_row_bitmap <= 16'b0000000000000000;
		15'h45ed: char_row_bitmap <= 16'b0000000000000000;
		15'h45ee: char_row_bitmap <= 16'b0000000000000000;
		15'h45ef: char_row_bitmap <= 16'b0000000000000000;
		15'h45f0: char_row_bitmap <= 16'b0000000000000000;
		15'h45f1: char_row_bitmap <= 16'b0000000000000000;
		15'h45f2: char_row_bitmap <= 16'b0000000000000000;
		15'h45f3: char_row_bitmap <= 16'b0000000000000000;
		15'h45f4: char_row_bitmap <= 16'b0000000000000000;
		15'h45f5: char_row_bitmap <= 16'b0000000000000000;
		15'h45f6: char_row_bitmap <= 16'b0000000000000000;
		15'h45f7: char_row_bitmap <= 16'b0000000000000000;
		15'h45f8: char_row_bitmap <= 16'b0000000000000000;
		15'h45f9: char_row_bitmap <= 16'b0000000000000000;
		15'h45fa: char_row_bitmap <= 16'b0000000000000000;
		15'h45fb: char_row_bitmap <= 16'b0000000000000000;
		15'h45fc: char_row_bitmap <= 16'b0000000000000000;
		15'h45fd: char_row_bitmap <= 16'b0000000000000000;
		15'h45fe: char_row_bitmap <= 16'b0000000000000000;
		15'h45ff: char_row_bitmap <= 16'b0000000000000000;
		15'h4600: char_row_bitmap <= 16'b0000000000000000;
		15'h4601: char_row_bitmap <= 16'b0000000000000000;
		15'h4602: char_row_bitmap <= 16'b0000000000000000;
		15'h4603: char_row_bitmap <= 16'b0000000000000000;
		15'h4604: char_row_bitmap <= 16'b0000000000000000;
		15'h4605: char_row_bitmap <= 16'b0000000000000000;
		15'h4606: char_row_bitmap <= 16'b0000000000000000;
		15'h4607: char_row_bitmap <= 16'b0000000000000000;
		15'h4608: char_row_bitmap <= 16'b0000000000000000;
		15'h4609: char_row_bitmap <= 16'b0000000000000000;
		15'h460a: char_row_bitmap <= 16'b0000000000000000;
		15'h460b: char_row_bitmap <= 16'b0000000000000000;
		15'h460c: char_row_bitmap <= 16'b0000000000000000;
		15'h460d: char_row_bitmap <= 16'b0000000000000000;
		15'h460e: char_row_bitmap <= 16'b0000000000000000;
		15'h460f: char_row_bitmap <= 16'b0000000000000000;
		15'h4610: char_row_bitmap <= 16'b0000000000000000;
		15'h4611: char_row_bitmap <= 16'b0000000000000000;
		15'h4612: char_row_bitmap <= 16'b0000000000000000;
		15'h4613: char_row_bitmap <= 16'b0000000000000000;
		15'h4614: char_row_bitmap <= 16'b0011111100000000;
		15'h4615: char_row_bitmap <= 16'b0011111100000000;
		15'h4616: char_row_bitmap <= 16'b0011111100000000;
		15'h4617: char_row_bitmap <= 16'b0011111100000000;
		15'h4618: char_row_bitmap <= 16'b0000000000000000;
		15'h4619: char_row_bitmap <= 16'b0000000000000000;
		15'h461a: char_row_bitmap <= 16'b0000000000000000;
		15'h461b: char_row_bitmap <= 16'b0000000000000000;
		15'h461c: char_row_bitmap <= 16'b0000000000000000;
		15'h461d: char_row_bitmap <= 16'b0000000000000000;
		15'h461e: char_row_bitmap <= 16'b0000000000000000;
		15'h461f: char_row_bitmap <= 16'b0000000000000000;
		15'h4620: char_row_bitmap <= 16'b0000000000000000;
		15'h4621: char_row_bitmap <= 16'b0000000000000000;
		15'h4622: char_row_bitmap <= 16'b0000000000000000;
		15'h4623: char_row_bitmap <= 16'b0000000000000000;
		15'h4624: char_row_bitmap <= 16'b0000000000000000;
		15'h4625: char_row_bitmap <= 16'b0000000000000000;
		15'h4626: char_row_bitmap <= 16'b0000000000000000;
		15'h4627: char_row_bitmap <= 16'b0000000000000000;
		15'h4628: char_row_bitmap <= 16'b0000000000111111;
		15'h4629: char_row_bitmap <= 16'b0000000000111111;
		15'h462a: char_row_bitmap <= 16'b0000000000111111;
		15'h462b: char_row_bitmap <= 16'b0000000000111111;
		15'h462c: char_row_bitmap <= 16'b0000000000000000;
		15'h462d: char_row_bitmap <= 16'b0000000000000000;
		15'h462e: char_row_bitmap <= 16'b0000000000000000;
		15'h462f: char_row_bitmap <= 16'b0000000000000000;
		15'h4630: char_row_bitmap <= 16'b0000000000000000;
		15'h4631: char_row_bitmap <= 16'b0000000000000000;
		15'h4632: char_row_bitmap <= 16'b0000000000000000;
		15'h4633: char_row_bitmap <= 16'b0000000000000000;
		15'h4634: char_row_bitmap <= 16'b0000000000000000;
		15'h4635: char_row_bitmap <= 16'b0000000000000000;
		15'h4636: char_row_bitmap <= 16'b0000000000000000;
		15'h4637: char_row_bitmap <= 16'b0000000000000000;
		15'h4638: char_row_bitmap <= 16'b0000000000000000;
		15'h4639: char_row_bitmap <= 16'b0000000000000000;
		15'h463a: char_row_bitmap <= 16'b0000000000000000;
		15'h463b: char_row_bitmap <= 16'b0000000000000000;
		15'h463c: char_row_bitmap <= 16'b0011111100111111;
		15'h463d: char_row_bitmap <= 16'b0011111100111111;
		15'h463e: char_row_bitmap <= 16'b0011111100111111;
		15'h463f: char_row_bitmap <= 16'b0011111100111111;
		15'h4640: char_row_bitmap <= 16'b0000000000000000;
		15'h4641: char_row_bitmap <= 16'b0000000000000000;
		15'h4642: char_row_bitmap <= 16'b0000000000000000;
		15'h4643: char_row_bitmap <= 16'b0000000000000000;
		15'h4644: char_row_bitmap <= 16'b0000000000000000;
		15'h4645: char_row_bitmap <= 16'b0000000000000000;
		15'h4646: char_row_bitmap <= 16'b0000000000000000;
		15'h4647: char_row_bitmap <= 16'b0000000000000000;
		15'h4648: char_row_bitmap <= 16'b0000000000000000;
		15'h4649: char_row_bitmap <= 16'b0000000000000000;
		15'h464a: char_row_bitmap <= 16'b0000000000000000;
		15'h464b: char_row_bitmap <= 16'b0000000000000000;
		15'h464c: char_row_bitmap <= 16'b0000000000000000;
		15'h464d: char_row_bitmap <= 16'b0000000000000000;
		15'h464e: char_row_bitmap <= 16'b0000000000000000;
		15'h464f: char_row_bitmap <= 16'b0000000000000000;
		15'h4650: char_row_bitmap <= 16'b0000000000000000;
		15'h4651: char_row_bitmap <= 16'b0000000000000000;
		15'h4652: char_row_bitmap <= 16'b0000000000000000;
		15'h4653: char_row_bitmap <= 16'b0000000000000000;
		15'h4654: char_row_bitmap <= 16'b0000000000000000;
		15'h4655: char_row_bitmap <= 16'b0000000000000000;
		15'h4656: char_row_bitmap <= 16'b0011111100000000;
		15'h4657: char_row_bitmap <= 16'b0011111100000000;
		15'h4658: char_row_bitmap <= 16'b0011111100000000;
		15'h4659: char_row_bitmap <= 16'b0011111100000000;
		15'h465a: char_row_bitmap <= 16'b0011111100000000;
		15'h465b: char_row_bitmap <= 16'b0011111100000000;
		15'h465c: char_row_bitmap <= 16'b0000000000000000;
		15'h465d: char_row_bitmap <= 16'b0000000000000000;
		15'h465e: char_row_bitmap <= 16'b0000000000000000;
		15'h465f: char_row_bitmap <= 16'b0000000000000000;
		15'h4660: char_row_bitmap <= 16'b0000000000000000;
		15'h4661: char_row_bitmap <= 16'b0000000000000000;
		15'h4662: char_row_bitmap <= 16'b0000000000000000;
		15'h4663: char_row_bitmap <= 16'b0000000000000000;
		15'h4664: char_row_bitmap <= 16'b0011111100000000;
		15'h4665: char_row_bitmap <= 16'b0011111100000000;
		15'h4666: char_row_bitmap <= 16'b0011111100000000;
		15'h4667: char_row_bitmap <= 16'b0011111100000000;
		15'h4668: char_row_bitmap <= 16'b0000000000000000;
		15'h4669: char_row_bitmap <= 16'b0000000000000000;
		15'h466a: char_row_bitmap <= 16'b0011111100000000;
		15'h466b: char_row_bitmap <= 16'b0011111100000000;
		15'h466c: char_row_bitmap <= 16'b0011111100000000;
		15'h466d: char_row_bitmap <= 16'b0011111100000000;
		15'h466e: char_row_bitmap <= 16'b0011111100000000;
		15'h466f: char_row_bitmap <= 16'b0011111100000000;
		15'h4670: char_row_bitmap <= 16'b0000000000000000;
		15'h4671: char_row_bitmap <= 16'b0000000000000000;
		15'h4672: char_row_bitmap <= 16'b0000000000000000;
		15'h4673: char_row_bitmap <= 16'b0000000000000000;
		15'h4674: char_row_bitmap <= 16'b0000000000000000;
		15'h4675: char_row_bitmap <= 16'b0000000000000000;
		15'h4676: char_row_bitmap <= 16'b0000000000000000;
		15'h4677: char_row_bitmap <= 16'b0000000000000000;
		15'h4678: char_row_bitmap <= 16'b0000000000111111;
		15'h4679: char_row_bitmap <= 16'b0000000000111111;
		15'h467a: char_row_bitmap <= 16'b0000000000111111;
		15'h467b: char_row_bitmap <= 16'b0000000000111111;
		15'h467c: char_row_bitmap <= 16'b0000000000000000;
		15'h467d: char_row_bitmap <= 16'b0000000000000000;
		15'h467e: char_row_bitmap <= 16'b0011111100000000;
		15'h467f: char_row_bitmap <= 16'b0011111100000000;
		15'h4680: char_row_bitmap <= 16'b0011111100000000;
		15'h4681: char_row_bitmap <= 16'b0011111100000000;
		15'h4682: char_row_bitmap <= 16'b0011111100000000;
		15'h4683: char_row_bitmap <= 16'b0011111100000000;
		15'h4684: char_row_bitmap <= 16'b0000000000000000;
		15'h4685: char_row_bitmap <= 16'b0000000000000000;
		15'h4686: char_row_bitmap <= 16'b0000000000000000;
		15'h4687: char_row_bitmap <= 16'b0000000000000000;
		15'h4688: char_row_bitmap <= 16'b0000000000000000;
		15'h4689: char_row_bitmap <= 16'b0000000000000000;
		15'h468a: char_row_bitmap <= 16'b0000000000000000;
		15'h468b: char_row_bitmap <= 16'b0000000000000000;
		15'h468c: char_row_bitmap <= 16'b0011111100111111;
		15'h468d: char_row_bitmap <= 16'b0011111100111111;
		15'h468e: char_row_bitmap <= 16'b0011111100111111;
		15'h468f: char_row_bitmap <= 16'b0011111100111111;
		15'h4690: char_row_bitmap <= 16'b0000000000000000;
		15'h4691: char_row_bitmap <= 16'b0000000000000000;
		15'h4692: char_row_bitmap <= 16'b0011111100000000;
		15'h4693: char_row_bitmap <= 16'b0011111100000000;
		15'h4694: char_row_bitmap <= 16'b0011111100000000;
		15'h4695: char_row_bitmap <= 16'b0011111100000000;
		15'h4696: char_row_bitmap <= 16'b0011111100000000;
		15'h4697: char_row_bitmap <= 16'b0011111100000000;
		15'h4698: char_row_bitmap <= 16'b0000000000000000;
		15'h4699: char_row_bitmap <= 16'b0000000000000000;
		15'h469a: char_row_bitmap <= 16'b0000000000000000;
		15'h469b: char_row_bitmap <= 16'b0000000000000000;
		15'h469c: char_row_bitmap <= 16'b0000000000000000;
		15'h469d: char_row_bitmap <= 16'b0000000000000000;
		15'h469e: char_row_bitmap <= 16'b0000000000000000;
		15'h469f: char_row_bitmap <= 16'b0000000000000000;
		15'h46a0: char_row_bitmap <= 16'b0000000000000000;
		15'h46a1: char_row_bitmap <= 16'b0000000000000000;
		15'h46a2: char_row_bitmap <= 16'b0000000000000000;
		15'h46a3: char_row_bitmap <= 16'b0000000000000000;
		15'h46a4: char_row_bitmap <= 16'b0000000000000000;
		15'h46a5: char_row_bitmap <= 16'b0000000000000000;
		15'h46a6: char_row_bitmap <= 16'b0000000000111111;
		15'h46a7: char_row_bitmap <= 16'b0000000000111111;
		15'h46a8: char_row_bitmap <= 16'b0000000000111111;
		15'h46a9: char_row_bitmap <= 16'b0000000000111111;
		15'h46aa: char_row_bitmap <= 16'b0000000000111111;
		15'h46ab: char_row_bitmap <= 16'b0000000000111111;
		15'h46ac: char_row_bitmap <= 16'b0000000000000000;
		15'h46ad: char_row_bitmap <= 16'b0000000000000000;
		15'h46ae: char_row_bitmap <= 16'b0000000000000000;
		15'h46af: char_row_bitmap <= 16'b0000000000000000;
		15'h46b0: char_row_bitmap <= 16'b0000000000000000;
		15'h46b1: char_row_bitmap <= 16'b0000000000000000;
		15'h46b2: char_row_bitmap <= 16'b0000000000000000;
		15'h46b3: char_row_bitmap <= 16'b0000000000000000;
		15'h46b4: char_row_bitmap <= 16'b0011111100000000;
		15'h46b5: char_row_bitmap <= 16'b0011111100000000;
		15'h46b6: char_row_bitmap <= 16'b0011111100000000;
		15'h46b7: char_row_bitmap <= 16'b0011111100000000;
		15'h46b8: char_row_bitmap <= 16'b0000000000000000;
		15'h46b9: char_row_bitmap <= 16'b0000000000000000;
		15'h46ba: char_row_bitmap <= 16'b0000000000111111;
		15'h46bb: char_row_bitmap <= 16'b0000000000111111;
		15'h46bc: char_row_bitmap <= 16'b0000000000111111;
		15'h46bd: char_row_bitmap <= 16'b0000000000111111;
		15'h46be: char_row_bitmap <= 16'b0000000000111111;
		15'h46bf: char_row_bitmap <= 16'b0000000000111111;
		15'h46c0: char_row_bitmap <= 16'b0000000000000000;
		15'h46c1: char_row_bitmap <= 16'b0000000000000000;
		15'h46c2: char_row_bitmap <= 16'b0000000000000000;
		15'h46c3: char_row_bitmap <= 16'b0000000000000000;
		15'h46c4: char_row_bitmap <= 16'b0000000000000000;
		15'h46c5: char_row_bitmap <= 16'b0000000000000000;
		15'h46c6: char_row_bitmap <= 16'b0000000000000000;
		15'h46c7: char_row_bitmap <= 16'b0000000000000000;
		15'h46c8: char_row_bitmap <= 16'b0000000000111111;
		15'h46c9: char_row_bitmap <= 16'b0000000000111111;
		15'h46ca: char_row_bitmap <= 16'b0000000000111111;
		15'h46cb: char_row_bitmap <= 16'b0000000000111111;
		15'h46cc: char_row_bitmap <= 16'b0000000000000000;
		15'h46cd: char_row_bitmap <= 16'b0000000000000000;
		15'h46ce: char_row_bitmap <= 16'b0000000000111111;
		15'h46cf: char_row_bitmap <= 16'b0000000000111111;
		15'h46d0: char_row_bitmap <= 16'b0000000000111111;
		15'h46d1: char_row_bitmap <= 16'b0000000000111111;
		15'h46d2: char_row_bitmap <= 16'b0000000000111111;
		15'h46d3: char_row_bitmap <= 16'b0000000000111111;
		15'h46d4: char_row_bitmap <= 16'b0000000000000000;
		15'h46d5: char_row_bitmap <= 16'b0000000000000000;
		15'h46d6: char_row_bitmap <= 16'b0000000000000000;
		15'h46d7: char_row_bitmap <= 16'b0000000000000000;
		15'h46d8: char_row_bitmap <= 16'b0000000000000000;
		15'h46d9: char_row_bitmap <= 16'b0000000000000000;
		15'h46da: char_row_bitmap <= 16'b0000000000000000;
		15'h46db: char_row_bitmap <= 16'b0000000000000000;
		15'h46dc: char_row_bitmap <= 16'b0011111100111111;
		15'h46dd: char_row_bitmap <= 16'b0011111100111111;
		15'h46de: char_row_bitmap <= 16'b0011111100111111;
		15'h46df: char_row_bitmap <= 16'b0011111100111111;
		15'h46e0: char_row_bitmap <= 16'b0000000000000000;
		15'h46e1: char_row_bitmap <= 16'b0000000000000000;
		15'h46e2: char_row_bitmap <= 16'b0000000000111111;
		15'h46e3: char_row_bitmap <= 16'b0000000000111111;
		15'h46e4: char_row_bitmap <= 16'b0000000000111111;
		15'h46e5: char_row_bitmap <= 16'b0000000000111111;
		15'h46e6: char_row_bitmap <= 16'b0000000000111111;
		15'h46e7: char_row_bitmap <= 16'b0000000000111111;
		15'h46e8: char_row_bitmap <= 16'b0000000000000000;
		15'h46e9: char_row_bitmap <= 16'b0000000000000000;
		15'h46ea: char_row_bitmap <= 16'b0000000000000000;
		15'h46eb: char_row_bitmap <= 16'b0000000000000000;
		15'h46ec: char_row_bitmap <= 16'b0000000000000000;
		15'h46ed: char_row_bitmap <= 16'b0000000000000000;
		15'h46ee: char_row_bitmap <= 16'b0000000000000000;
		15'h46ef: char_row_bitmap <= 16'b0000000000000000;
		15'h46f0: char_row_bitmap <= 16'b0000000000000000;
		15'h46f1: char_row_bitmap <= 16'b0000000000000000;
		15'h46f2: char_row_bitmap <= 16'b0000000000000000;
		15'h46f3: char_row_bitmap <= 16'b0000000000000000;
		15'h46f4: char_row_bitmap <= 16'b0000000000000000;
		15'h46f5: char_row_bitmap <= 16'b0000000000000000;
		15'h46f6: char_row_bitmap <= 16'b0011111100111111;
		15'h46f7: char_row_bitmap <= 16'b0011111100111111;
		15'h46f8: char_row_bitmap <= 16'b0011111100111111;
		15'h46f9: char_row_bitmap <= 16'b0011111100111111;
		15'h46fa: char_row_bitmap <= 16'b0011111100111111;
		15'h46fb: char_row_bitmap <= 16'b0011111100111111;
		15'h46fc: char_row_bitmap <= 16'b0000000000000000;
		15'h46fd: char_row_bitmap <= 16'b0000000000000000;
		15'h46fe: char_row_bitmap <= 16'b0000000000000000;
		15'h46ff: char_row_bitmap <= 16'b0000000000000000;
		15'h4700: char_row_bitmap <= 16'b0000000000000000;
		15'h4701: char_row_bitmap <= 16'b0000000000000000;
		15'h4702: char_row_bitmap <= 16'b0000000000000000;
		15'h4703: char_row_bitmap <= 16'b0000000000000000;
		15'h4704: char_row_bitmap <= 16'b0011111100000000;
		15'h4705: char_row_bitmap <= 16'b0011111100000000;
		15'h4706: char_row_bitmap <= 16'b0011111100000000;
		15'h4707: char_row_bitmap <= 16'b0011111100000000;
		15'h4708: char_row_bitmap <= 16'b0000000000000000;
		15'h4709: char_row_bitmap <= 16'b0000000000000000;
		15'h470a: char_row_bitmap <= 16'b0011111100111111;
		15'h470b: char_row_bitmap <= 16'b0011111100111111;
		15'h470c: char_row_bitmap <= 16'b0011111100111111;
		15'h470d: char_row_bitmap <= 16'b0011111100111111;
		15'h470e: char_row_bitmap <= 16'b0011111100111111;
		15'h470f: char_row_bitmap <= 16'b0011111100111111;
		15'h4710: char_row_bitmap <= 16'b0000000000000000;
		15'h4711: char_row_bitmap <= 16'b0000000000000000;
		15'h4712: char_row_bitmap <= 16'b0000000000000000;
		15'h4713: char_row_bitmap <= 16'b0000000000000000;
		15'h4714: char_row_bitmap <= 16'b0000000000000000;
		15'h4715: char_row_bitmap <= 16'b0000000000000000;
		15'h4716: char_row_bitmap <= 16'b0000000000000000;
		15'h4717: char_row_bitmap <= 16'b0000000000000000;
		15'h4718: char_row_bitmap <= 16'b0000000000111111;
		15'h4719: char_row_bitmap <= 16'b0000000000111111;
		15'h471a: char_row_bitmap <= 16'b0000000000111111;
		15'h471b: char_row_bitmap <= 16'b0000000000111111;
		15'h471c: char_row_bitmap <= 16'b0000000000000000;
		15'h471d: char_row_bitmap <= 16'b0000000000000000;
		15'h471e: char_row_bitmap <= 16'b0011111100111111;
		15'h471f: char_row_bitmap <= 16'b0011111100111111;
		15'h4720: char_row_bitmap <= 16'b0011111100111111;
		15'h4721: char_row_bitmap <= 16'b0011111100111111;
		15'h4722: char_row_bitmap <= 16'b0011111100111111;
		15'h4723: char_row_bitmap <= 16'b0011111100111111;
		15'h4724: char_row_bitmap <= 16'b0000000000000000;
		15'h4725: char_row_bitmap <= 16'b0000000000000000;
		15'h4726: char_row_bitmap <= 16'b0000000000000000;
		15'h4727: char_row_bitmap <= 16'b0000000000000000;
		15'h4728: char_row_bitmap <= 16'b0000000000000000;
		15'h4729: char_row_bitmap <= 16'b0000000000000000;
		15'h472a: char_row_bitmap <= 16'b0000000000000000;
		15'h472b: char_row_bitmap <= 16'b0000000000000000;
		15'h472c: char_row_bitmap <= 16'b0011111100111111;
		15'h472d: char_row_bitmap <= 16'b0011111100111111;
		15'h472e: char_row_bitmap <= 16'b0011111100111111;
		15'h472f: char_row_bitmap <= 16'b0011111100111111;
		15'h4730: char_row_bitmap <= 16'b0000000000000000;
		15'h4731: char_row_bitmap <= 16'b0000000000000000;
		15'h4732: char_row_bitmap <= 16'b0011111100111111;
		15'h4733: char_row_bitmap <= 16'b0011111100111111;
		15'h4734: char_row_bitmap <= 16'b0011111100111111;
		15'h4735: char_row_bitmap <= 16'b0011111100111111;
		15'h4736: char_row_bitmap <= 16'b0011111100111111;
		15'h4737: char_row_bitmap <= 16'b0011111100111111;
		15'h4738: char_row_bitmap <= 16'b0000000000000000;
		15'h4739: char_row_bitmap <= 16'b0000000000000000;
		15'h473a: char_row_bitmap <= 16'b0000000000000000;
		15'h473b: char_row_bitmap <= 16'b0000000000000000;
		15'h473c: char_row_bitmap <= 16'b0000000000000000;
		15'h473d: char_row_bitmap <= 16'b0000000000000000;
		15'h473e: char_row_bitmap <= 16'b0000000000000000;
		15'h473f: char_row_bitmap <= 16'b0000000000000000;
		15'h4740: char_row_bitmap <= 16'b0000000000000000;
		15'h4741: char_row_bitmap <= 16'b0000000000000000;
		15'h4742: char_row_bitmap <= 16'b0000000000000000;
		15'h4743: char_row_bitmap <= 16'b0000000000000000;
		15'h4744: char_row_bitmap <= 16'b0000000000000000;
		15'h4745: char_row_bitmap <= 16'b0000000000000000;
		15'h4746: char_row_bitmap <= 16'b0000000000000000;
		15'h4747: char_row_bitmap <= 16'b0000000000000000;
		15'h4748: char_row_bitmap <= 16'b0000000000000000;
		15'h4749: char_row_bitmap <= 16'b0000000000000000;
		15'h474a: char_row_bitmap <= 16'b0000000000000000;
		15'h474b: char_row_bitmap <= 16'b0000000000000000;
		15'h474c: char_row_bitmap <= 16'b0000000000000000;
		15'h474d: char_row_bitmap <= 16'b0000000000000000;
		15'h474e: char_row_bitmap <= 16'b0011111100000000;
		15'h474f: char_row_bitmap <= 16'b0011111100000000;
		15'h4750: char_row_bitmap <= 16'b0011111100000000;
		15'h4751: char_row_bitmap <= 16'b0011111100000000;
		15'h4752: char_row_bitmap <= 16'b0000000000000000;
		15'h4753: char_row_bitmap <= 16'b0000000000000000;
		15'h4754: char_row_bitmap <= 16'b0011111100000000;
		15'h4755: char_row_bitmap <= 16'b0011111100000000;
		15'h4756: char_row_bitmap <= 16'b0011111100000000;
		15'h4757: char_row_bitmap <= 16'b0011111100000000;
		15'h4758: char_row_bitmap <= 16'b0000000000000000;
		15'h4759: char_row_bitmap <= 16'b0000000000000000;
		15'h475a: char_row_bitmap <= 16'b0000000000000000;
		15'h475b: char_row_bitmap <= 16'b0000000000000000;
		15'h475c: char_row_bitmap <= 16'b0000000000000000;
		15'h475d: char_row_bitmap <= 16'b0000000000000000;
		15'h475e: char_row_bitmap <= 16'b0000000000000000;
		15'h475f: char_row_bitmap <= 16'b0000000000000000;
		15'h4760: char_row_bitmap <= 16'b0000000000000000;
		15'h4761: char_row_bitmap <= 16'b0000000000000000;
		15'h4762: char_row_bitmap <= 16'b0011111100000000;
		15'h4763: char_row_bitmap <= 16'b0011111100000000;
		15'h4764: char_row_bitmap <= 16'b0011111100000000;
		15'h4765: char_row_bitmap <= 16'b0011111100000000;
		15'h4766: char_row_bitmap <= 16'b0000000000000000;
		15'h4767: char_row_bitmap <= 16'b0000000000000000;
		15'h4768: char_row_bitmap <= 16'b0000000000111111;
		15'h4769: char_row_bitmap <= 16'b0000000000111111;
		15'h476a: char_row_bitmap <= 16'b0000000000111111;
		15'h476b: char_row_bitmap <= 16'b0000000000111111;
		15'h476c: char_row_bitmap <= 16'b0000000000000000;
		15'h476d: char_row_bitmap <= 16'b0000000000000000;
		15'h476e: char_row_bitmap <= 16'b0000000000000000;
		15'h476f: char_row_bitmap <= 16'b0000000000000000;
		15'h4770: char_row_bitmap <= 16'b0000000000000000;
		15'h4771: char_row_bitmap <= 16'b0000000000000000;
		15'h4772: char_row_bitmap <= 16'b0000000000000000;
		15'h4773: char_row_bitmap <= 16'b0000000000000000;
		15'h4774: char_row_bitmap <= 16'b0000000000000000;
		15'h4775: char_row_bitmap <= 16'b0000000000000000;
		15'h4776: char_row_bitmap <= 16'b0011111100000000;
		15'h4777: char_row_bitmap <= 16'b0011111100000000;
		15'h4778: char_row_bitmap <= 16'b0011111100000000;
		15'h4779: char_row_bitmap <= 16'b0011111100000000;
		15'h477a: char_row_bitmap <= 16'b0000000000000000;
		15'h477b: char_row_bitmap <= 16'b0000000000000000;
		15'h477c: char_row_bitmap <= 16'b0011111100111111;
		15'h477d: char_row_bitmap <= 16'b0011111100111111;
		15'h477e: char_row_bitmap <= 16'b0011111100111111;
		15'h477f: char_row_bitmap <= 16'b0011111100111111;
		15'h4780: char_row_bitmap <= 16'b0000000000000000;
		15'h4781: char_row_bitmap <= 16'b0000000000000000;
		15'h4782: char_row_bitmap <= 16'b0000000000000000;
		15'h4783: char_row_bitmap <= 16'b0000000000000000;
		15'h4784: char_row_bitmap <= 16'b0000000000000000;
		15'h4785: char_row_bitmap <= 16'b0000000000000000;
		15'h4786: char_row_bitmap <= 16'b0000000000000000;
		15'h4787: char_row_bitmap <= 16'b0000000000000000;
		15'h4788: char_row_bitmap <= 16'b0000000000000000;
		15'h4789: char_row_bitmap <= 16'b0000000000000000;
		15'h478a: char_row_bitmap <= 16'b0011111100000000;
		15'h478b: char_row_bitmap <= 16'b0011111100000000;
		15'h478c: char_row_bitmap <= 16'b0011111100000000;
		15'h478d: char_row_bitmap <= 16'b0011111100000000;
		15'h478e: char_row_bitmap <= 16'b0000000000000000;
		15'h478f: char_row_bitmap <= 16'b0000000000000000;
		15'h4790: char_row_bitmap <= 16'b0000000000000000;
		15'h4791: char_row_bitmap <= 16'b0000000000000000;
		15'h4792: char_row_bitmap <= 16'b0000000000000000;
		15'h4793: char_row_bitmap <= 16'b0000000000000000;
		15'h4794: char_row_bitmap <= 16'b0000000000000000;
		15'h4795: char_row_bitmap <= 16'b0000000000000000;
		15'h4796: char_row_bitmap <= 16'b0011111100000000;
		15'h4797: char_row_bitmap <= 16'b0011111100000000;
		15'h4798: char_row_bitmap <= 16'b0011111100000000;
		15'h4799: char_row_bitmap <= 16'b0011111100000000;
		15'h479a: char_row_bitmap <= 16'b0011111100000000;
		15'h479b: char_row_bitmap <= 16'b0011111100000000;
		15'h479c: char_row_bitmap <= 16'b0000000000000000;
		15'h479d: char_row_bitmap <= 16'b0000000000000000;
		15'h479e: char_row_bitmap <= 16'b0011111100000000;
		15'h479f: char_row_bitmap <= 16'b0011111100000000;
		15'h47a0: char_row_bitmap <= 16'b0011111100000000;
		15'h47a1: char_row_bitmap <= 16'b0011111100000000;
		15'h47a2: char_row_bitmap <= 16'b0000000000000000;
		15'h47a3: char_row_bitmap <= 16'b0000000000000000;
		15'h47a4: char_row_bitmap <= 16'b0011111100000000;
		15'h47a5: char_row_bitmap <= 16'b0011111100000000;
		15'h47a6: char_row_bitmap <= 16'b0011111100000000;
		15'h47a7: char_row_bitmap <= 16'b0011111100000000;
		15'h47a8: char_row_bitmap <= 16'b0000000000000000;
		15'h47a9: char_row_bitmap <= 16'b0000000000000000;
		15'h47aa: char_row_bitmap <= 16'b0011111100000000;
		15'h47ab: char_row_bitmap <= 16'b0011111100000000;
		15'h47ac: char_row_bitmap <= 16'b0011111100000000;
		15'h47ad: char_row_bitmap <= 16'b0011111100000000;
		15'h47ae: char_row_bitmap <= 16'b0011111100000000;
		15'h47af: char_row_bitmap <= 16'b0011111100000000;
		15'h47b0: char_row_bitmap <= 16'b0000000000000000;
		15'h47b1: char_row_bitmap <= 16'b0000000000000000;
		15'h47b2: char_row_bitmap <= 16'b0011111100000000;
		15'h47b3: char_row_bitmap <= 16'b0011111100000000;
		15'h47b4: char_row_bitmap <= 16'b0011111100000000;
		15'h47b5: char_row_bitmap <= 16'b0011111100000000;
		15'h47b6: char_row_bitmap <= 16'b0000000000000000;
		15'h47b7: char_row_bitmap <= 16'b0000000000000000;
		15'h47b8: char_row_bitmap <= 16'b0000000000111111;
		15'h47b9: char_row_bitmap <= 16'b0000000000111111;
		15'h47ba: char_row_bitmap <= 16'b0000000000111111;
		15'h47bb: char_row_bitmap <= 16'b0000000000111111;
		15'h47bc: char_row_bitmap <= 16'b0000000000000000;
		15'h47bd: char_row_bitmap <= 16'b0000000000000000;
		15'h47be: char_row_bitmap <= 16'b0011111100000000;
		15'h47bf: char_row_bitmap <= 16'b0011111100000000;
		15'h47c0: char_row_bitmap <= 16'b0011111100000000;
		15'h47c1: char_row_bitmap <= 16'b0011111100000000;
		15'h47c2: char_row_bitmap <= 16'b0011111100000000;
		15'h47c3: char_row_bitmap <= 16'b0011111100000000;
		15'h47c4: char_row_bitmap <= 16'b0000000000000000;
		15'h47c5: char_row_bitmap <= 16'b0000000000000000;
		15'h47c6: char_row_bitmap <= 16'b0011111100000000;
		15'h47c7: char_row_bitmap <= 16'b0011111100000000;
		15'h47c8: char_row_bitmap <= 16'b0011111100000000;
		15'h47c9: char_row_bitmap <= 16'b0011111100000000;
		15'h47ca: char_row_bitmap <= 16'b0000000000000000;
		15'h47cb: char_row_bitmap <= 16'b0000000000000000;
		15'h47cc: char_row_bitmap <= 16'b0011111100111111;
		15'h47cd: char_row_bitmap <= 16'b0011111100111111;
		15'h47ce: char_row_bitmap <= 16'b0011111100111111;
		15'h47cf: char_row_bitmap <= 16'b0011111100111111;
		15'h47d0: char_row_bitmap <= 16'b0000000000000000;
		15'h47d1: char_row_bitmap <= 16'b0000000000000000;
		15'h47d2: char_row_bitmap <= 16'b0011111100000000;
		15'h47d3: char_row_bitmap <= 16'b0011111100000000;
		15'h47d4: char_row_bitmap <= 16'b0011111100000000;
		15'h47d5: char_row_bitmap <= 16'b0011111100000000;
		15'h47d6: char_row_bitmap <= 16'b0011111100000000;
		15'h47d7: char_row_bitmap <= 16'b0011111100000000;
		15'h47d8: char_row_bitmap <= 16'b0000000000000000;
		15'h47d9: char_row_bitmap <= 16'b0000000000000000;
		15'h47da: char_row_bitmap <= 16'b0011111100000000;
		15'h47db: char_row_bitmap <= 16'b0011111100000000;
		15'h47dc: char_row_bitmap <= 16'b0011111100000000;
		15'h47dd: char_row_bitmap <= 16'b0011111100000000;
		15'h47de: char_row_bitmap <= 16'b0000000000000000;
		15'h47df: char_row_bitmap <= 16'b0000000000000000;
		15'h47e0: char_row_bitmap <= 16'b0000000000000000;
		15'h47e1: char_row_bitmap <= 16'b0000000000000000;
		15'h47e2: char_row_bitmap <= 16'b0000000000000000;
		15'h47e3: char_row_bitmap <= 16'b0000000000000000;
		15'h47e4: char_row_bitmap <= 16'b0000000000000000;
		15'h47e5: char_row_bitmap <= 16'b0000000000000000;
		15'h47e6: char_row_bitmap <= 16'b0000000000111111;
		15'h47e7: char_row_bitmap <= 16'b0000000000111111;
		15'h47e8: char_row_bitmap <= 16'b0000000000111111;
		15'h47e9: char_row_bitmap <= 16'b0000000000111111;
		15'h47ea: char_row_bitmap <= 16'b0000000000111111;
		15'h47eb: char_row_bitmap <= 16'b0000000000111111;
		15'h47ec: char_row_bitmap <= 16'b0000000000000000;
		15'h47ed: char_row_bitmap <= 16'b0000000000000000;
		15'h47ee: char_row_bitmap <= 16'b0011111100000000;
		15'h47ef: char_row_bitmap <= 16'b0011111100000000;
		15'h47f0: char_row_bitmap <= 16'b0011111100000000;
		15'h47f1: char_row_bitmap <= 16'b0011111100000000;
		15'h47f2: char_row_bitmap <= 16'b0000000000000000;
		15'h47f3: char_row_bitmap <= 16'b0000000000000000;
		15'h47f4: char_row_bitmap <= 16'b0011111100000000;
		15'h47f5: char_row_bitmap <= 16'b0011111100000000;
		15'h47f6: char_row_bitmap <= 16'b0011111100000000;
		15'h47f7: char_row_bitmap <= 16'b0011111100000000;
		15'h47f8: char_row_bitmap <= 16'b0000000000000000;
		15'h47f9: char_row_bitmap <= 16'b0000000000000000;
		15'h47fa: char_row_bitmap <= 16'b0000000000111111;
		15'h47fb: char_row_bitmap <= 16'b0000000000111111;
		15'h47fc: char_row_bitmap <= 16'b0000000000111111;
		15'h47fd: char_row_bitmap <= 16'b0000000000111111;
		15'h47fe: char_row_bitmap <= 16'b0000000000111111;
		15'h47ff: char_row_bitmap <= 16'b0000000000111111;
		15'h4800: char_row_bitmap <= 16'b0000000000000000;
		15'h4801: char_row_bitmap <= 16'b0000000000000000;
		15'h4802: char_row_bitmap <= 16'b0011111100000000;
		15'h4803: char_row_bitmap <= 16'b0011111100000000;
		15'h4804: char_row_bitmap <= 16'b0011111100000000;
		15'h4805: char_row_bitmap <= 16'b0011111100000000;
		15'h4806: char_row_bitmap <= 16'b0000000000000000;
		15'h4807: char_row_bitmap <= 16'b0000000000000000;
		15'h4808: char_row_bitmap <= 16'b0000000000111111;
		15'h4809: char_row_bitmap <= 16'b0000000000111111;
		15'h480a: char_row_bitmap <= 16'b0000000000111111;
		15'h480b: char_row_bitmap <= 16'b0000000000111111;
		15'h480c: char_row_bitmap <= 16'b0000000000000000;
		15'h480d: char_row_bitmap <= 16'b0000000000000000;
		15'h480e: char_row_bitmap <= 16'b0000000000111111;
		15'h480f: char_row_bitmap <= 16'b0000000000111111;
		15'h4810: char_row_bitmap <= 16'b0000000000111111;
		15'h4811: char_row_bitmap <= 16'b0000000000111111;
		15'h4812: char_row_bitmap <= 16'b0000000000111111;
		15'h4813: char_row_bitmap <= 16'b0000000000111111;
		15'h4814: char_row_bitmap <= 16'b0000000000000000;
		15'h4815: char_row_bitmap <= 16'b0000000000000000;
		15'h4816: char_row_bitmap <= 16'b0011111100000000;
		15'h4817: char_row_bitmap <= 16'b0011111100000000;
		15'h4818: char_row_bitmap <= 16'b0011111100000000;
		15'h4819: char_row_bitmap <= 16'b0011111100000000;
		15'h481a: char_row_bitmap <= 16'b0000000000000000;
		15'h481b: char_row_bitmap <= 16'b0000000000000000;
		15'h481c: char_row_bitmap <= 16'b0011111100111111;
		15'h481d: char_row_bitmap <= 16'b0011111100111111;
		15'h481e: char_row_bitmap <= 16'b0011111100111111;
		15'h481f: char_row_bitmap <= 16'b0011111100111111;
		15'h4820: char_row_bitmap <= 16'b0000000000000000;
		15'h4821: char_row_bitmap <= 16'b0000000000000000;
		15'h4822: char_row_bitmap <= 16'b0000000000111111;
		15'h4823: char_row_bitmap <= 16'b0000000000111111;
		15'h4824: char_row_bitmap <= 16'b0000000000111111;
		15'h4825: char_row_bitmap <= 16'b0000000000111111;
		15'h4826: char_row_bitmap <= 16'b0000000000111111;
		15'h4827: char_row_bitmap <= 16'b0000000000111111;
		15'h4828: char_row_bitmap <= 16'b0000000000000000;
		15'h4829: char_row_bitmap <= 16'b0000000000000000;
		15'h482a: char_row_bitmap <= 16'b0011111100000000;
		15'h482b: char_row_bitmap <= 16'b0011111100000000;
		15'h482c: char_row_bitmap <= 16'b0011111100000000;
		15'h482d: char_row_bitmap <= 16'b0011111100000000;
		15'h482e: char_row_bitmap <= 16'b0000000000000000;
		15'h482f: char_row_bitmap <= 16'b0000000000000000;
		15'h4830: char_row_bitmap <= 16'b0000000000000000;
		15'h4831: char_row_bitmap <= 16'b0000000000000000;
		15'h4832: char_row_bitmap <= 16'b0000000000000000;
		15'h4833: char_row_bitmap <= 16'b0000000000000000;
		15'h4834: char_row_bitmap <= 16'b0000000000000000;
		15'h4835: char_row_bitmap <= 16'b0000000000000000;
		15'h4836: char_row_bitmap <= 16'b0011111100111111;
		15'h4837: char_row_bitmap <= 16'b0011111100111111;
		15'h4838: char_row_bitmap <= 16'b0011111100111111;
		15'h4839: char_row_bitmap <= 16'b0011111100111111;
		15'h483a: char_row_bitmap <= 16'b0011111100111111;
		15'h483b: char_row_bitmap <= 16'b0011111100111111;
		15'h483c: char_row_bitmap <= 16'b0000000000000000;
		15'h483d: char_row_bitmap <= 16'b0000000000000000;
		15'h483e: char_row_bitmap <= 16'b0011111100000000;
		15'h483f: char_row_bitmap <= 16'b0011111100000000;
		15'h4840: char_row_bitmap <= 16'b0011111100000000;
		15'h4841: char_row_bitmap <= 16'b0011111100000000;
		15'h4842: char_row_bitmap <= 16'b0000000000000000;
		15'h4843: char_row_bitmap <= 16'b0000000000000000;
		15'h4844: char_row_bitmap <= 16'b0011111100000000;
		15'h4845: char_row_bitmap <= 16'b0011111100000000;
		15'h4846: char_row_bitmap <= 16'b0011111100000000;
		15'h4847: char_row_bitmap <= 16'b0011111100000000;
		15'h4848: char_row_bitmap <= 16'b0000000000000000;
		15'h4849: char_row_bitmap <= 16'b0000000000000000;
		15'h484a: char_row_bitmap <= 16'b0011111100111111;
		15'h484b: char_row_bitmap <= 16'b0011111100111111;
		15'h484c: char_row_bitmap <= 16'b0011111100111111;
		15'h484d: char_row_bitmap <= 16'b0011111100111111;
		15'h484e: char_row_bitmap <= 16'b0011111100111111;
		15'h484f: char_row_bitmap <= 16'b0011111100111111;
		15'h4850: char_row_bitmap <= 16'b0000000000000000;
		15'h4851: char_row_bitmap <= 16'b0000000000000000;
		15'h4852: char_row_bitmap <= 16'b0011111100000000;
		15'h4853: char_row_bitmap <= 16'b0011111100000000;
		15'h4854: char_row_bitmap <= 16'b0011111100000000;
		15'h4855: char_row_bitmap <= 16'b0011111100000000;
		15'h4856: char_row_bitmap <= 16'b0000000000000000;
		15'h4857: char_row_bitmap <= 16'b0000000000000000;
		15'h4858: char_row_bitmap <= 16'b0000000000111111;
		15'h4859: char_row_bitmap <= 16'b0000000000111111;
		15'h485a: char_row_bitmap <= 16'b0000000000111111;
		15'h485b: char_row_bitmap <= 16'b0000000000111111;
		15'h485c: char_row_bitmap <= 16'b0000000000000000;
		15'h485d: char_row_bitmap <= 16'b0000000000000000;
		15'h485e: char_row_bitmap <= 16'b0011111100111111;
		15'h485f: char_row_bitmap <= 16'b0011111100111111;
		15'h4860: char_row_bitmap <= 16'b0011111100111111;
		15'h4861: char_row_bitmap <= 16'b0011111100111111;
		15'h4862: char_row_bitmap <= 16'b0011111100111111;
		15'h4863: char_row_bitmap <= 16'b0011111100111111;
		15'h4864: char_row_bitmap <= 16'b0000000000000000;
		15'h4865: char_row_bitmap <= 16'b0000000000000000;
		15'h4866: char_row_bitmap <= 16'b0011111100000000;
		15'h4867: char_row_bitmap <= 16'b0011111100000000;
		15'h4868: char_row_bitmap <= 16'b0011111100000000;
		15'h4869: char_row_bitmap <= 16'b0011111100000000;
		15'h486a: char_row_bitmap <= 16'b0000000000000000;
		15'h486b: char_row_bitmap <= 16'b0000000000000000;
		15'h486c: char_row_bitmap <= 16'b0011111100111111;
		15'h486d: char_row_bitmap <= 16'b0011111100111111;
		15'h486e: char_row_bitmap <= 16'b0011111100111111;
		15'h486f: char_row_bitmap <= 16'b0011111100111111;
		15'h4870: char_row_bitmap <= 16'b0000000000000000;
		15'h4871: char_row_bitmap <= 16'b0000000000000000;
		15'h4872: char_row_bitmap <= 16'b0011111100111111;
		15'h4873: char_row_bitmap <= 16'b0011111100111111;
		15'h4874: char_row_bitmap <= 16'b0011111100111111;
		15'h4875: char_row_bitmap <= 16'b0011111100111111;
		15'h4876: char_row_bitmap <= 16'b0011111100111111;
		15'h4877: char_row_bitmap <= 16'b0011111100111111;
		15'h4878: char_row_bitmap <= 16'b0000000000000000;
		15'h4879: char_row_bitmap <= 16'b0000000000000000;
		15'h487a: char_row_bitmap <= 16'b0011111100000000;
		15'h487b: char_row_bitmap <= 16'b0011111100000000;
		15'h487c: char_row_bitmap <= 16'b0011111100000000;
		15'h487d: char_row_bitmap <= 16'b0011111100000000;
		15'h487e: char_row_bitmap <= 16'b0000000000000000;
		15'h487f: char_row_bitmap <= 16'b0000000000000000;
		15'h4880: char_row_bitmap <= 16'b0000000000000000;
		15'h4881: char_row_bitmap <= 16'b0000000000000000;
		15'h4882: char_row_bitmap <= 16'b0000000000000000;
		15'h4883: char_row_bitmap <= 16'b0000000000000000;
		15'h4884: char_row_bitmap <= 16'b0000000000000000;
		15'h4885: char_row_bitmap <= 16'b0000000000000000;
		15'h4886: char_row_bitmap <= 16'b0000000000000000;
		15'h4887: char_row_bitmap <= 16'b0000000000000000;
		15'h4888: char_row_bitmap <= 16'b0000000000000000;
		15'h4889: char_row_bitmap <= 16'b0000000000000000;
		15'h488a: char_row_bitmap <= 16'b0000000000000000;
		15'h488b: char_row_bitmap <= 16'b0000000000000000;
		15'h488c: char_row_bitmap <= 16'b0000000000000000;
		15'h488d: char_row_bitmap <= 16'b0000000000000000;
		15'h488e: char_row_bitmap <= 16'b0000000000111111;
		15'h488f: char_row_bitmap <= 16'b0000000000111111;
		15'h4890: char_row_bitmap <= 16'b0000000000111111;
		15'h4891: char_row_bitmap <= 16'b0000000000111111;
		15'h4892: char_row_bitmap <= 16'b0000000000000000;
		15'h4893: char_row_bitmap <= 16'b0000000000000000;
		15'h4894: char_row_bitmap <= 16'b0011111100000000;
		15'h4895: char_row_bitmap <= 16'b0011111100000000;
		15'h4896: char_row_bitmap <= 16'b0011111100000000;
		15'h4897: char_row_bitmap <= 16'b0011111100000000;
		15'h4898: char_row_bitmap <= 16'b0000000000000000;
		15'h4899: char_row_bitmap <= 16'b0000000000000000;
		15'h489a: char_row_bitmap <= 16'b0000000000000000;
		15'h489b: char_row_bitmap <= 16'b0000000000000000;
		15'h489c: char_row_bitmap <= 16'b0000000000000000;
		15'h489d: char_row_bitmap <= 16'b0000000000000000;
		15'h489e: char_row_bitmap <= 16'b0000000000000000;
		15'h489f: char_row_bitmap <= 16'b0000000000000000;
		15'h48a0: char_row_bitmap <= 16'b0000000000000000;
		15'h48a1: char_row_bitmap <= 16'b0000000000000000;
		15'h48a2: char_row_bitmap <= 16'b0000000000111111;
		15'h48a3: char_row_bitmap <= 16'b0000000000111111;
		15'h48a4: char_row_bitmap <= 16'b0000000000111111;
		15'h48a5: char_row_bitmap <= 16'b0000000000111111;
		15'h48a6: char_row_bitmap <= 16'b0000000000000000;
		15'h48a7: char_row_bitmap <= 16'b0000000000000000;
		15'h48a8: char_row_bitmap <= 16'b0000000000111111;
		15'h48a9: char_row_bitmap <= 16'b0000000000111111;
		15'h48aa: char_row_bitmap <= 16'b0000000000111111;
		15'h48ab: char_row_bitmap <= 16'b0000000000111111;
		15'h48ac: char_row_bitmap <= 16'b0000000000000000;
		15'h48ad: char_row_bitmap <= 16'b0000000000000000;
		15'h48ae: char_row_bitmap <= 16'b0000000000000000;
		15'h48af: char_row_bitmap <= 16'b0000000000000000;
		15'h48b0: char_row_bitmap <= 16'b0000000000000000;
		15'h48b1: char_row_bitmap <= 16'b0000000000000000;
		15'h48b2: char_row_bitmap <= 16'b0000000000000000;
		15'h48b3: char_row_bitmap <= 16'b0000000000000000;
		15'h48b4: char_row_bitmap <= 16'b0000000000000000;
		15'h48b5: char_row_bitmap <= 16'b0000000000000000;
		15'h48b6: char_row_bitmap <= 16'b0000000000111111;
		15'h48b7: char_row_bitmap <= 16'b0000000000111111;
		15'h48b8: char_row_bitmap <= 16'b0000000000111111;
		15'h48b9: char_row_bitmap <= 16'b0000000000111111;
		15'h48ba: char_row_bitmap <= 16'b0000000000000000;
		15'h48bb: char_row_bitmap <= 16'b0000000000000000;
		15'h48bc: char_row_bitmap <= 16'b0011111100111111;
		15'h48bd: char_row_bitmap <= 16'b0011111100111111;
		15'h48be: char_row_bitmap <= 16'b0011111100111111;
		15'h48bf: char_row_bitmap <= 16'b0011111100111111;
		15'h48c0: char_row_bitmap <= 16'b0000000000000000;
		15'h48c1: char_row_bitmap <= 16'b0000000000000000;
		15'h48c2: char_row_bitmap <= 16'b0000000000000000;
		15'h48c3: char_row_bitmap <= 16'b0000000000000000;
		15'h48c4: char_row_bitmap <= 16'b0000000000000000;
		15'h48c5: char_row_bitmap <= 16'b0000000000000000;
		15'h48c6: char_row_bitmap <= 16'b0000000000000000;
		15'h48c7: char_row_bitmap <= 16'b0000000000000000;
		15'h48c8: char_row_bitmap <= 16'b0000000000000000;
		15'h48c9: char_row_bitmap <= 16'b0000000000000000;
		15'h48ca: char_row_bitmap <= 16'b0000000000111111;
		15'h48cb: char_row_bitmap <= 16'b0000000000111111;
		15'h48cc: char_row_bitmap <= 16'b0000000000111111;
		15'h48cd: char_row_bitmap <= 16'b0000000000111111;
		15'h48ce: char_row_bitmap <= 16'b0000000000000000;
		15'h48cf: char_row_bitmap <= 16'b0000000000000000;
		15'h48d0: char_row_bitmap <= 16'b0000000000000000;
		15'h48d1: char_row_bitmap <= 16'b0000000000000000;
		15'h48d2: char_row_bitmap <= 16'b0000000000000000;
		15'h48d3: char_row_bitmap <= 16'b0000000000000000;
		15'h48d4: char_row_bitmap <= 16'b0000000000000000;
		15'h48d5: char_row_bitmap <= 16'b0000000000000000;
		15'h48d6: char_row_bitmap <= 16'b0011111100000000;
		15'h48d7: char_row_bitmap <= 16'b0011111100000000;
		15'h48d8: char_row_bitmap <= 16'b0011111100000000;
		15'h48d9: char_row_bitmap <= 16'b0011111100000000;
		15'h48da: char_row_bitmap <= 16'b0011111100000000;
		15'h48db: char_row_bitmap <= 16'b0011111100000000;
		15'h48dc: char_row_bitmap <= 16'b0000000000000000;
		15'h48dd: char_row_bitmap <= 16'b0000000000000000;
		15'h48de: char_row_bitmap <= 16'b0000000000111111;
		15'h48df: char_row_bitmap <= 16'b0000000000111111;
		15'h48e0: char_row_bitmap <= 16'b0000000000111111;
		15'h48e1: char_row_bitmap <= 16'b0000000000111111;
		15'h48e2: char_row_bitmap <= 16'b0000000000000000;
		15'h48e3: char_row_bitmap <= 16'b0000000000000000;
		15'h48e4: char_row_bitmap <= 16'b0011111100000000;
		15'h48e5: char_row_bitmap <= 16'b0011111100000000;
		15'h48e6: char_row_bitmap <= 16'b0011111100000000;
		15'h48e7: char_row_bitmap <= 16'b0011111100000000;
		15'h48e8: char_row_bitmap <= 16'b0000000000000000;
		15'h48e9: char_row_bitmap <= 16'b0000000000000000;
		15'h48ea: char_row_bitmap <= 16'b0011111100000000;
		15'h48eb: char_row_bitmap <= 16'b0011111100000000;
		15'h48ec: char_row_bitmap <= 16'b0011111100000000;
		15'h48ed: char_row_bitmap <= 16'b0011111100000000;
		15'h48ee: char_row_bitmap <= 16'b0011111100000000;
		15'h48ef: char_row_bitmap <= 16'b0011111100000000;
		15'h48f0: char_row_bitmap <= 16'b0000000000000000;
		15'h48f1: char_row_bitmap <= 16'b0000000000000000;
		15'h48f2: char_row_bitmap <= 16'b0000000000111111;
		15'h48f3: char_row_bitmap <= 16'b0000000000111111;
		15'h48f4: char_row_bitmap <= 16'b0000000000111111;
		15'h48f5: char_row_bitmap <= 16'b0000000000111111;
		15'h48f6: char_row_bitmap <= 16'b0000000000000000;
		15'h48f7: char_row_bitmap <= 16'b0000000000000000;
		15'h48f8: char_row_bitmap <= 16'b0000000000111111;
		15'h48f9: char_row_bitmap <= 16'b0000000000111111;
		15'h48fa: char_row_bitmap <= 16'b0000000000111111;
		15'h48fb: char_row_bitmap <= 16'b0000000000111111;
		15'h48fc: char_row_bitmap <= 16'b0000000000000000;
		15'h48fd: char_row_bitmap <= 16'b0000000000000000;
		15'h48fe: char_row_bitmap <= 16'b0011111100000000;
		15'h48ff: char_row_bitmap <= 16'b0011111100000000;
		15'h4900: char_row_bitmap <= 16'b0011111100000000;
		15'h4901: char_row_bitmap <= 16'b0011111100000000;
		15'h4902: char_row_bitmap <= 16'b0011111100000000;
		15'h4903: char_row_bitmap <= 16'b0011111100000000;
		15'h4904: char_row_bitmap <= 16'b0000000000000000;
		15'h4905: char_row_bitmap <= 16'b0000000000000000;
		15'h4906: char_row_bitmap <= 16'b0000000000111111;
		15'h4907: char_row_bitmap <= 16'b0000000000111111;
		15'h4908: char_row_bitmap <= 16'b0000000000111111;
		15'h4909: char_row_bitmap <= 16'b0000000000111111;
		15'h490a: char_row_bitmap <= 16'b0000000000000000;
		15'h490b: char_row_bitmap <= 16'b0000000000000000;
		15'h490c: char_row_bitmap <= 16'b0011111100111111;
		15'h490d: char_row_bitmap <= 16'b0011111100111111;
		15'h490e: char_row_bitmap <= 16'b0011111100111111;
		15'h490f: char_row_bitmap <= 16'b0011111100111111;
		15'h4910: char_row_bitmap <= 16'b0000000000000000;
		15'h4911: char_row_bitmap <= 16'b0000000000000000;
		15'h4912: char_row_bitmap <= 16'b0011111100000000;
		15'h4913: char_row_bitmap <= 16'b0011111100000000;
		15'h4914: char_row_bitmap <= 16'b0011111100000000;
		15'h4915: char_row_bitmap <= 16'b0011111100000000;
		15'h4916: char_row_bitmap <= 16'b0011111100000000;
		15'h4917: char_row_bitmap <= 16'b0011111100000000;
		15'h4918: char_row_bitmap <= 16'b0000000000000000;
		15'h4919: char_row_bitmap <= 16'b0000000000000000;
		15'h491a: char_row_bitmap <= 16'b0000000000111111;
		15'h491b: char_row_bitmap <= 16'b0000000000111111;
		15'h491c: char_row_bitmap <= 16'b0000000000111111;
		15'h491d: char_row_bitmap <= 16'b0000000000111111;
		15'h491e: char_row_bitmap <= 16'b0000000000000000;
		15'h491f: char_row_bitmap <= 16'b0000000000000000;
		15'h4920: char_row_bitmap <= 16'b0000000000000000;
		15'h4921: char_row_bitmap <= 16'b0000000000000000;
		15'h4922: char_row_bitmap <= 16'b0000000000000000;
		15'h4923: char_row_bitmap <= 16'b0000000000000000;
		15'h4924: char_row_bitmap <= 16'b0000000000000000;
		15'h4925: char_row_bitmap <= 16'b0000000000000000;
		15'h4926: char_row_bitmap <= 16'b0000000000111111;
		15'h4927: char_row_bitmap <= 16'b0000000000111111;
		15'h4928: char_row_bitmap <= 16'b0000000000111111;
		15'h4929: char_row_bitmap <= 16'b0000000000111111;
		15'h492a: char_row_bitmap <= 16'b0000000000111111;
		15'h492b: char_row_bitmap <= 16'b0000000000111111;
		15'h492c: char_row_bitmap <= 16'b0000000000000000;
		15'h492d: char_row_bitmap <= 16'b0000000000000000;
		15'h492e: char_row_bitmap <= 16'b0000000000111111;
		15'h492f: char_row_bitmap <= 16'b0000000000111111;
		15'h4930: char_row_bitmap <= 16'b0000000000111111;
		15'h4931: char_row_bitmap <= 16'b0000000000111111;
		15'h4932: char_row_bitmap <= 16'b0000000000000000;
		15'h4933: char_row_bitmap <= 16'b0000000000000000;
		15'h4934: char_row_bitmap <= 16'b0011111100000000;
		15'h4935: char_row_bitmap <= 16'b0011111100000000;
		15'h4936: char_row_bitmap <= 16'b0011111100000000;
		15'h4937: char_row_bitmap <= 16'b0011111100000000;
		15'h4938: char_row_bitmap <= 16'b0000000000000000;
		15'h4939: char_row_bitmap <= 16'b0000000000000000;
		15'h493a: char_row_bitmap <= 16'b0000000000111111;
		15'h493b: char_row_bitmap <= 16'b0000000000111111;
		15'h493c: char_row_bitmap <= 16'b0000000000111111;
		15'h493d: char_row_bitmap <= 16'b0000000000111111;
		15'h493e: char_row_bitmap <= 16'b0000000000111111;
		15'h493f: char_row_bitmap <= 16'b0000000000111111;
		15'h4940: char_row_bitmap <= 16'b0000000000000000;
		15'h4941: char_row_bitmap <= 16'b0000000000000000;
		15'h4942: char_row_bitmap <= 16'b0000000000111111;
		15'h4943: char_row_bitmap <= 16'b0000000000111111;
		15'h4944: char_row_bitmap <= 16'b0000000000111111;
		15'h4945: char_row_bitmap <= 16'b0000000000111111;
		15'h4946: char_row_bitmap <= 16'b0000000000000000;
		15'h4947: char_row_bitmap <= 16'b0000000000000000;
		15'h4948: char_row_bitmap <= 16'b0000000000111111;
		15'h4949: char_row_bitmap <= 16'b0000000000111111;
		15'h494a: char_row_bitmap <= 16'b0000000000111111;
		15'h494b: char_row_bitmap <= 16'b0000000000111111;
		15'h494c: char_row_bitmap <= 16'b0000000000000000;
		15'h494d: char_row_bitmap <= 16'b0000000000000000;
		15'h494e: char_row_bitmap <= 16'b0000000000111111;
		15'h494f: char_row_bitmap <= 16'b0000000000111111;
		15'h4950: char_row_bitmap <= 16'b0000000000111111;
		15'h4951: char_row_bitmap <= 16'b0000000000111111;
		15'h4952: char_row_bitmap <= 16'b0000000000111111;
		15'h4953: char_row_bitmap <= 16'b0000000000111111;
		15'h4954: char_row_bitmap <= 16'b0000000000000000;
		15'h4955: char_row_bitmap <= 16'b0000000000000000;
		15'h4956: char_row_bitmap <= 16'b0000000000111111;
		15'h4957: char_row_bitmap <= 16'b0000000000111111;
		15'h4958: char_row_bitmap <= 16'b0000000000111111;
		15'h4959: char_row_bitmap <= 16'b0000000000111111;
		15'h495a: char_row_bitmap <= 16'b0000000000000000;
		15'h495b: char_row_bitmap <= 16'b0000000000000000;
		15'h495c: char_row_bitmap <= 16'b0011111100111111;
		15'h495d: char_row_bitmap <= 16'b0011111100111111;
		15'h495e: char_row_bitmap <= 16'b0011111100111111;
		15'h495f: char_row_bitmap <= 16'b0011111100111111;
		15'h4960: char_row_bitmap <= 16'b0000000000000000;
		15'h4961: char_row_bitmap <= 16'b0000000000000000;
		15'h4962: char_row_bitmap <= 16'b0000000000111111;
		15'h4963: char_row_bitmap <= 16'b0000000000111111;
		15'h4964: char_row_bitmap <= 16'b0000000000111111;
		15'h4965: char_row_bitmap <= 16'b0000000000111111;
		15'h4966: char_row_bitmap <= 16'b0000000000111111;
		15'h4967: char_row_bitmap <= 16'b0000000000111111;
		15'h4968: char_row_bitmap <= 16'b0000000000000000;
		15'h4969: char_row_bitmap <= 16'b0000000000000000;
		15'h496a: char_row_bitmap <= 16'b0000000000111111;
		15'h496b: char_row_bitmap <= 16'b0000000000111111;
		15'h496c: char_row_bitmap <= 16'b0000000000111111;
		15'h496d: char_row_bitmap <= 16'b0000000000111111;
		15'h496e: char_row_bitmap <= 16'b0000000000000000;
		15'h496f: char_row_bitmap <= 16'b0000000000000000;
		15'h4970: char_row_bitmap <= 16'b0000000000000000;
		15'h4971: char_row_bitmap <= 16'b0000000000000000;
		15'h4972: char_row_bitmap <= 16'b0000000000000000;
		15'h4973: char_row_bitmap <= 16'b0000000000000000;
		15'h4974: char_row_bitmap <= 16'b0000000000000000;
		15'h4975: char_row_bitmap <= 16'b0000000000000000;
		15'h4976: char_row_bitmap <= 16'b0011111100111111;
		15'h4977: char_row_bitmap <= 16'b0011111100111111;
		15'h4978: char_row_bitmap <= 16'b0011111100111111;
		15'h4979: char_row_bitmap <= 16'b0011111100111111;
		15'h497a: char_row_bitmap <= 16'b0011111100111111;
		15'h497b: char_row_bitmap <= 16'b0011111100111111;
		15'h497c: char_row_bitmap <= 16'b0000000000000000;
		15'h497d: char_row_bitmap <= 16'b0000000000000000;
		15'h497e: char_row_bitmap <= 16'b0000000000111111;
		15'h497f: char_row_bitmap <= 16'b0000000000111111;
		15'h4980: char_row_bitmap <= 16'b0000000000111111;
		15'h4981: char_row_bitmap <= 16'b0000000000111111;
		15'h4982: char_row_bitmap <= 16'b0000000000000000;
		15'h4983: char_row_bitmap <= 16'b0000000000000000;
		15'h4984: char_row_bitmap <= 16'b0011111100000000;
		15'h4985: char_row_bitmap <= 16'b0011111100000000;
		15'h4986: char_row_bitmap <= 16'b0011111100000000;
		15'h4987: char_row_bitmap <= 16'b0011111100000000;
		15'h4988: char_row_bitmap <= 16'b0000000000000000;
		15'h4989: char_row_bitmap <= 16'b0000000000000000;
		15'h498a: char_row_bitmap <= 16'b0011111100111111;
		15'h498b: char_row_bitmap <= 16'b0011111100111111;
		15'h498c: char_row_bitmap <= 16'b0011111100111111;
		15'h498d: char_row_bitmap <= 16'b0011111100111111;
		15'h498e: char_row_bitmap <= 16'b0011111100111111;
		15'h498f: char_row_bitmap <= 16'b0011111100111111;
		15'h4990: char_row_bitmap <= 16'b0000000000000000;
		15'h4991: char_row_bitmap <= 16'b0000000000000000;
		15'h4992: char_row_bitmap <= 16'b0000000000111111;
		15'h4993: char_row_bitmap <= 16'b0000000000111111;
		15'h4994: char_row_bitmap <= 16'b0000000000111111;
		15'h4995: char_row_bitmap <= 16'b0000000000111111;
		15'h4996: char_row_bitmap <= 16'b0000000000000000;
		15'h4997: char_row_bitmap <= 16'b0000000000000000;
		15'h4998: char_row_bitmap <= 16'b0000000000111111;
		15'h4999: char_row_bitmap <= 16'b0000000000111111;
		15'h499a: char_row_bitmap <= 16'b0000000000111111;
		15'h499b: char_row_bitmap <= 16'b0000000000111111;
		15'h499c: char_row_bitmap <= 16'b0000000000000000;
		15'h499d: char_row_bitmap <= 16'b0000000000000000;
		15'h499e: char_row_bitmap <= 16'b0011111100111111;
		15'h499f: char_row_bitmap <= 16'b0011111100111111;
		15'h49a0: char_row_bitmap <= 16'b0011111100111111;
		15'h49a1: char_row_bitmap <= 16'b0011111100111111;
		15'h49a2: char_row_bitmap <= 16'b0011111100111111;
		15'h49a3: char_row_bitmap <= 16'b0011111100111111;
		15'h49a4: char_row_bitmap <= 16'b0000000000000000;
		15'h49a5: char_row_bitmap <= 16'b0000000000000000;
		15'h49a6: char_row_bitmap <= 16'b0000000000111111;
		15'h49a7: char_row_bitmap <= 16'b0000000000111111;
		15'h49a8: char_row_bitmap <= 16'b0000000000111111;
		15'h49a9: char_row_bitmap <= 16'b0000000000111111;
		15'h49aa: char_row_bitmap <= 16'b0000000000000000;
		15'h49ab: char_row_bitmap <= 16'b0000000000000000;
		15'h49ac: char_row_bitmap <= 16'b0011111100111111;
		15'h49ad: char_row_bitmap <= 16'b0011111100111111;
		15'h49ae: char_row_bitmap <= 16'b0011111100111111;
		15'h49af: char_row_bitmap <= 16'b0011111100111111;
		15'h49b0: char_row_bitmap <= 16'b0000000000000000;
		15'h49b1: char_row_bitmap <= 16'b0000000000000000;
		15'h49b2: char_row_bitmap <= 16'b0011111100111111;
		15'h49b3: char_row_bitmap <= 16'b0011111100111111;
		15'h49b4: char_row_bitmap <= 16'b0011111100111111;
		15'h49b5: char_row_bitmap <= 16'b0011111100111111;
		15'h49b6: char_row_bitmap <= 16'b0011111100111111;
		15'h49b7: char_row_bitmap <= 16'b0011111100111111;
		15'h49b8: char_row_bitmap <= 16'b0000000000000000;
		15'h49b9: char_row_bitmap <= 16'b0000000000000000;
		15'h49ba: char_row_bitmap <= 16'b0000000000111111;
		15'h49bb: char_row_bitmap <= 16'b0000000000111111;
		15'h49bc: char_row_bitmap <= 16'b0000000000111111;
		15'h49bd: char_row_bitmap <= 16'b0000000000111111;
		15'h49be: char_row_bitmap <= 16'b0000000000000000;
		15'h49bf: char_row_bitmap <= 16'b0000000000000000;
		15'h49c0: char_row_bitmap <= 16'b0000000000000000;
		15'h49c1: char_row_bitmap <= 16'b0000000000000000;
		15'h49c2: char_row_bitmap <= 16'b0000000000000000;
		15'h49c3: char_row_bitmap <= 16'b0000000000000000;
		15'h49c4: char_row_bitmap <= 16'b0000000000000000;
		15'h49c5: char_row_bitmap <= 16'b0000000000000000;
		15'h49c6: char_row_bitmap <= 16'b0000000000000000;
		15'h49c7: char_row_bitmap <= 16'b0000000000000000;
		15'h49c8: char_row_bitmap <= 16'b0000000000000000;
		15'h49c9: char_row_bitmap <= 16'b0000000000000000;
		15'h49ca: char_row_bitmap <= 16'b0000000000000000;
		15'h49cb: char_row_bitmap <= 16'b0000000000000000;
		15'h49cc: char_row_bitmap <= 16'b0000000000000000;
		15'h49cd: char_row_bitmap <= 16'b0000000000000000;
		15'h49ce: char_row_bitmap <= 16'b0011111100111111;
		15'h49cf: char_row_bitmap <= 16'b0011111100111111;
		15'h49d0: char_row_bitmap <= 16'b0011111100111111;
		15'h49d1: char_row_bitmap <= 16'b0011111100111111;
		15'h49d2: char_row_bitmap <= 16'b0000000000000000;
		15'h49d3: char_row_bitmap <= 16'b0000000000000000;
		15'h49d4: char_row_bitmap <= 16'b0011111100000000;
		15'h49d5: char_row_bitmap <= 16'b0011111100000000;
		15'h49d6: char_row_bitmap <= 16'b0011111100000000;
		15'h49d7: char_row_bitmap <= 16'b0011111100000000;
		15'h49d8: char_row_bitmap <= 16'b0000000000000000;
		15'h49d9: char_row_bitmap <= 16'b0000000000000000;
		15'h49da: char_row_bitmap <= 16'b0000000000000000;
		15'h49db: char_row_bitmap <= 16'b0000000000000000;
		15'h49dc: char_row_bitmap <= 16'b0000000000000000;
		15'h49dd: char_row_bitmap <= 16'b0000000000000000;
		15'h49de: char_row_bitmap <= 16'b0000000000000000;
		15'h49df: char_row_bitmap <= 16'b0000000000000000;
		15'h49e0: char_row_bitmap <= 16'b0000000000000000;
		15'h49e1: char_row_bitmap <= 16'b0000000000000000;
		15'h49e2: char_row_bitmap <= 16'b0011111100111111;
		15'h49e3: char_row_bitmap <= 16'b0011111100111111;
		15'h49e4: char_row_bitmap <= 16'b0011111100111111;
		15'h49e5: char_row_bitmap <= 16'b0011111100111111;
		15'h49e6: char_row_bitmap <= 16'b0000000000000000;
		15'h49e7: char_row_bitmap <= 16'b0000000000000000;
		15'h49e8: char_row_bitmap <= 16'b0000000000111111;
		15'h49e9: char_row_bitmap <= 16'b0000000000111111;
		15'h49ea: char_row_bitmap <= 16'b0000000000111111;
		15'h49eb: char_row_bitmap <= 16'b0000000000111111;
		15'h49ec: char_row_bitmap <= 16'b0000000000000000;
		15'h49ed: char_row_bitmap <= 16'b0000000000000000;
		15'h49ee: char_row_bitmap <= 16'b0000000000000000;
		15'h49ef: char_row_bitmap <= 16'b0000000000000000;
		15'h49f0: char_row_bitmap <= 16'b0000000000000000;
		15'h49f1: char_row_bitmap <= 16'b0000000000000000;
		15'h49f2: char_row_bitmap <= 16'b0000000000000000;
		15'h49f3: char_row_bitmap <= 16'b0000000000000000;
		15'h49f4: char_row_bitmap <= 16'b0000000000000000;
		15'h49f5: char_row_bitmap <= 16'b0000000000000000;
		15'h49f6: char_row_bitmap <= 16'b0011111100111111;
		15'h49f7: char_row_bitmap <= 16'b0011111100111111;
		15'h49f8: char_row_bitmap <= 16'b0011111100111111;
		15'h49f9: char_row_bitmap <= 16'b0011111100111111;
		15'h49fa: char_row_bitmap <= 16'b0000000000000000;
		15'h49fb: char_row_bitmap <= 16'b0000000000000000;
		15'h49fc: char_row_bitmap <= 16'b0011111100111111;
		15'h49fd: char_row_bitmap <= 16'b0011111100111111;
		15'h49fe: char_row_bitmap <= 16'b0011111100111111;
		15'h49ff: char_row_bitmap <= 16'b0011111100111111;
		15'h4a00: char_row_bitmap <= 16'b0000000000000000;
		15'h4a01: char_row_bitmap <= 16'b0000000000000000;
		15'h4a02: char_row_bitmap <= 16'b0000000000000000;
		15'h4a03: char_row_bitmap <= 16'b0000000000000000;
		15'h4a04: char_row_bitmap <= 16'b0000000000000000;
		15'h4a05: char_row_bitmap <= 16'b0000000000000000;
		15'h4a06: char_row_bitmap <= 16'b0000000000000000;
		15'h4a07: char_row_bitmap <= 16'b0000000000000000;
		15'h4a08: char_row_bitmap <= 16'b0000000000000000;
		15'h4a09: char_row_bitmap <= 16'b0000000000000000;
		15'h4a0a: char_row_bitmap <= 16'b0011111100111111;
		15'h4a0b: char_row_bitmap <= 16'b0011111100111111;
		15'h4a0c: char_row_bitmap <= 16'b0011111100111111;
		15'h4a0d: char_row_bitmap <= 16'b0011111100111111;
		15'h4a0e: char_row_bitmap <= 16'b0000000000000000;
		15'h4a0f: char_row_bitmap <= 16'b0000000000000000;
		15'h4a10: char_row_bitmap <= 16'b0000000000000000;
		15'h4a11: char_row_bitmap <= 16'b0000000000000000;
		15'h4a12: char_row_bitmap <= 16'b0000000000000000;
		15'h4a13: char_row_bitmap <= 16'b0000000000000000;
		15'h4a14: char_row_bitmap <= 16'b0000000000000000;
		15'h4a15: char_row_bitmap <= 16'b0000000000000000;
		15'h4a16: char_row_bitmap <= 16'b0011111100000000;
		15'h4a17: char_row_bitmap <= 16'b0011111100000000;
		15'h4a18: char_row_bitmap <= 16'b0011111100000000;
		15'h4a19: char_row_bitmap <= 16'b0011111100000000;
		15'h4a1a: char_row_bitmap <= 16'b0011111100000000;
		15'h4a1b: char_row_bitmap <= 16'b0011111100000000;
		15'h4a1c: char_row_bitmap <= 16'b0000000000000000;
		15'h4a1d: char_row_bitmap <= 16'b0000000000000000;
		15'h4a1e: char_row_bitmap <= 16'b0011111100111111;
		15'h4a1f: char_row_bitmap <= 16'b0011111100111111;
		15'h4a20: char_row_bitmap <= 16'b0011111100111111;
		15'h4a21: char_row_bitmap <= 16'b0011111100111111;
		15'h4a22: char_row_bitmap <= 16'b0000000000000000;
		15'h4a23: char_row_bitmap <= 16'b0000000000000000;
		15'h4a24: char_row_bitmap <= 16'b0011111100000000;
		15'h4a25: char_row_bitmap <= 16'b0011111100000000;
		15'h4a26: char_row_bitmap <= 16'b0011111100000000;
		15'h4a27: char_row_bitmap <= 16'b0011111100000000;
		15'h4a28: char_row_bitmap <= 16'b0000000000000000;
		15'h4a29: char_row_bitmap <= 16'b0000000000000000;
		15'h4a2a: char_row_bitmap <= 16'b0011111100000000;
		15'h4a2b: char_row_bitmap <= 16'b0011111100000000;
		15'h4a2c: char_row_bitmap <= 16'b0011111100000000;
		15'h4a2d: char_row_bitmap <= 16'b0011111100000000;
		15'h4a2e: char_row_bitmap <= 16'b0011111100000000;
		15'h4a2f: char_row_bitmap <= 16'b0011111100000000;
		15'h4a30: char_row_bitmap <= 16'b0000000000000000;
		15'h4a31: char_row_bitmap <= 16'b0000000000000000;
		15'h4a32: char_row_bitmap <= 16'b0011111100111111;
		15'h4a33: char_row_bitmap <= 16'b0011111100111111;
		15'h4a34: char_row_bitmap <= 16'b0011111100111111;
		15'h4a35: char_row_bitmap <= 16'b0011111100111111;
		15'h4a36: char_row_bitmap <= 16'b0000000000000000;
		15'h4a37: char_row_bitmap <= 16'b0000000000000000;
		15'h4a38: char_row_bitmap <= 16'b0000000000111111;
		15'h4a39: char_row_bitmap <= 16'b0000000000111111;
		15'h4a3a: char_row_bitmap <= 16'b0000000000111111;
		15'h4a3b: char_row_bitmap <= 16'b0000000000111111;
		15'h4a3c: char_row_bitmap <= 16'b0000000000000000;
		15'h4a3d: char_row_bitmap <= 16'b0000000000000000;
		15'h4a3e: char_row_bitmap <= 16'b0011111100000000;
		15'h4a3f: char_row_bitmap <= 16'b0011111100000000;
		15'h4a40: char_row_bitmap <= 16'b0011111100000000;
		15'h4a41: char_row_bitmap <= 16'b0011111100000000;
		15'h4a42: char_row_bitmap <= 16'b0011111100000000;
		15'h4a43: char_row_bitmap <= 16'b0011111100000000;
		15'h4a44: char_row_bitmap <= 16'b0000000000000000;
		15'h4a45: char_row_bitmap <= 16'b0000000000000000;
		15'h4a46: char_row_bitmap <= 16'b0011111100111111;
		15'h4a47: char_row_bitmap <= 16'b0011111100111111;
		15'h4a48: char_row_bitmap <= 16'b0011111100111111;
		15'h4a49: char_row_bitmap <= 16'b0011111100111111;
		15'h4a4a: char_row_bitmap <= 16'b0000000000000000;
		15'h4a4b: char_row_bitmap <= 16'b0000000000000000;
		15'h4a4c: char_row_bitmap <= 16'b0011111100111111;
		15'h4a4d: char_row_bitmap <= 16'b0011111100111111;
		15'h4a4e: char_row_bitmap <= 16'b0011111100111111;
		15'h4a4f: char_row_bitmap <= 16'b0011111100111111;
		15'h4a50: char_row_bitmap <= 16'b0000000000000000;
		15'h4a51: char_row_bitmap <= 16'b0000000000000000;
		15'h4a52: char_row_bitmap <= 16'b0011111100000000;
		15'h4a53: char_row_bitmap <= 16'b0011111100000000;
		15'h4a54: char_row_bitmap <= 16'b0011111100000000;
		15'h4a55: char_row_bitmap <= 16'b0011111100000000;
		15'h4a56: char_row_bitmap <= 16'b0011111100000000;
		15'h4a57: char_row_bitmap <= 16'b0011111100000000;
		15'h4a58: char_row_bitmap <= 16'b0000000000000000;
		15'h4a59: char_row_bitmap <= 16'b0000000000000000;
		15'h4a5a: char_row_bitmap <= 16'b0011111100111111;
		15'h4a5b: char_row_bitmap <= 16'b0011111100111111;
		15'h4a5c: char_row_bitmap <= 16'b0011111100111111;
		15'h4a5d: char_row_bitmap <= 16'b0011111100111111;
		15'h4a5e: char_row_bitmap <= 16'b0000000000000000;
		15'h4a5f: char_row_bitmap <= 16'b0000000000000000;
		15'h4a60: char_row_bitmap <= 16'b0000000000000000;
		15'h4a61: char_row_bitmap <= 16'b0000000000000000;
		15'h4a62: char_row_bitmap <= 16'b0000000000000000;
		15'h4a63: char_row_bitmap <= 16'b0000000000000000;
		15'h4a64: char_row_bitmap <= 16'b0000000000000000;
		15'h4a65: char_row_bitmap <= 16'b0000000000000000;
		15'h4a66: char_row_bitmap <= 16'b0000000000111111;
		15'h4a67: char_row_bitmap <= 16'b0000000000111111;
		15'h4a68: char_row_bitmap <= 16'b0000000000111111;
		15'h4a69: char_row_bitmap <= 16'b0000000000111111;
		15'h4a6a: char_row_bitmap <= 16'b0000000000111111;
		15'h4a6b: char_row_bitmap <= 16'b0000000000111111;
		15'h4a6c: char_row_bitmap <= 16'b0000000000000000;
		15'h4a6d: char_row_bitmap <= 16'b0000000000000000;
		15'h4a6e: char_row_bitmap <= 16'b0011111100111111;
		15'h4a6f: char_row_bitmap <= 16'b0011111100111111;
		15'h4a70: char_row_bitmap <= 16'b0011111100111111;
		15'h4a71: char_row_bitmap <= 16'b0011111100111111;
		15'h4a72: char_row_bitmap <= 16'b0000000000000000;
		15'h4a73: char_row_bitmap <= 16'b0000000000000000;
		15'h4a74: char_row_bitmap <= 16'b0011111100000000;
		15'h4a75: char_row_bitmap <= 16'b0011111100000000;
		15'h4a76: char_row_bitmap <= 16'b0011111100000000;
		15'h4a77: char_row_bitmap <= 16'b0011111100000000;
		15'h4a78: char_row_bitmap <= 16'b0000000000000000;
		15'h4a79: char_row_bitmap <= 16'b0000000000000000;
		15'h4a7a: char_row_bitmap <= 16'b0000000000111111;
		15'h4a7b: char_row_bitmap <= 16'b0000000000111111;
		15'h4a7c: char_row_bitmap <= 16'b0000000000111111;
		15'h4a7d: char_row_bitmap <= 16'b0000000000111111;
		15'h4a7e: char_row_bitmap <= 16'b0000000000111111;
		15'h4a7f: char_row_bitmap <= 16'b0000000000111111;
		15'h4a80: char_row_bitmap <= 16'b0000000000000000;
		15'h4a81: char_row_bitmap <= 16'b0000000000000000;
		15'h4a82: char_row_bitmap <= 16'b0011111100111111;
		15'h4a83: char_row_bitmap <= 16'b0011111100111111;
		15'h4a84: char_row_bitmap <= 16'b0011111100111111;
		15'h4a85: char_row_bitmap <= 16'b0011111100111111;
		15'h4a86: char_row_bitmap <= 16'b0000000000000000;
		15'h4a87: char_row_bitmap <= 16'b0000000000000000;
		15'h4a88: char_row_bitmap <= 16'b0000000000111111;
		15'h4a89: char_row_bitmap <= 16'b0000000000111111;
		15'h4a8a: char_row_bitmap <= 16'b0000000000111111;
		15'h4a8b: char_row_bitmap <= 16'b0000000000111111;
		15'h4a8c: char_row_bitmap <= 16'b0000000000000000;
		15'h4a8d: char_row_bitmap <= 16'b0000000000000000;
		15'h4a8e: char_row_bitmap <= 16'b0000000000111111;
		15'h4a8f: char_row_bitmap <= 16'b0000000000111111;
		15'h4a90: char_row_bitmap <= 16'b0000000000111111;
		15'h4a91: char_row_bitmap <= 16'b0000000000111111;
		15'h4a92: char_row_bitmap <= 16'b0000000000111111;
		15'h4a93: char_row_bitmap <= 16'b0000000000111111;
		15'h4a94: char_row_bitmap <= 16'b0000000000000000;
		15'h4a95: char_row_bitmap <= 16'b0000000000000000;
		15'h4a96: char_row_bitmap <= 16'b0011111100111111;
		15'h4a97: char_row_bitmap <= 16'b0011111100111111;
		15'h4a98: char_row_bitmap <= 16'b0011111100111111;
		15'h4a99: char_row_bitmap <= 16'b0011111100111111;
		15'h4a9a: char_row_bitmap <= 16'b0000000000000000;
		15'h4a9b: char_row_bitmap <= 16'b0000000000000000;
		15'h4a9c: char_row_bitmap <= 16'b0011111100111111;
		15'h4a9d: char_row_bitmap <= 16'b0011111100111111;
		15'h4a9e: char_row_bitmap <= 16'b0011111100111111;
		15'h4a9f: char_row_bitmap <= 16'b0011111100111111;
		15'h4aa0: char_row_bitmap <= 16'b0000000000000000;
		15'h4aa1: char_row_bitmap <= 16'b0000000000000000;
		15'h4aa2: char_row_bitmap <= 16'b0000000000111111;
		15'h4aa3: char_row_bitmap <= 16'b0000000000111111;
		15'h4aa4: char_row_bitmap <= 16'b0000000000111111;
		15'h4aa5: char_row_bitmap <= 16'b0000000000111111;
		15'h4aa6: char_row_bitmap <= 16'b0000000000111111;
		15'h4aa7: char_row_bitmap <= 16'b0000000000111111;
		15'h4aa8: char_row_bitmap <= 16'b0000000000000000;
		15'h4aa9: char_row_bitmap <= 16'b0000000000000000;
		15'h4aaa: char_row_bitmap <= 16'b0011111100111111;
		15'h4aab: char_row_bitmap <= 16'b0011111100111111;
		15'h4aac: char_row_bitmap <= 16'b0011111100111111;
		15'h4aad: char_row_bitmap <= 16'b0011111100111111;
		15'h4aae: char_row_bitmap <= 16'b0000000000000000;
		15'h4aaf: char_row_bitmap <= 16'b0000000000000000;
		15'h4ab0: char_row_bitmap <= 16'b0000000000000000;
		15'h4ab1: char_row_bitmap <= 16'b0000000000000000;
		15'h4ab2: char_row_bitmap <= 16'b0000000000000000;
		15'h4ab3: char_row_bitmap <= 16'b0000000000000000;
		15'h4ab4: char_row_bitmap <= 16'b0000000000000000;
		15'h4ab5: char_row_bitmap <= 16'b0000000000000000;
		15'h4ab6: char_row_bitmap <= 16'b0011111100111111;
		15'h4ab7: char_row_bitmap <= 16'b0011111100111111;
		15'h4ab8: char_row_bitmap <= 16'b0011111100111111;
		15'h4ab9: char_row_bitmap <= 16'b0011111100111111;
		15'h4aba: char_row_bitmap <= 16'b0011111100111111;
		15'h4abb: char_row_bitmap <= 16'b0011111100111111;
		15'h4abc: char_row_bitmap <= 16'b0000000000000000;
		15'h4abd: char_row_bitmap <= 16'b0000000000000000;
		15'h4abe: char_row_bitmap <= 16'b0011111100111111;
		15'h4abf: char_row_bitmap <= 16'b0011111100111111;
		15'h4ac0: char_row_bitmap <= 16'b0011111100111111;
		15'h4ac1: char_row_bitmap <= 16'b0011111100111111;
		15'h4ac2: char_row_bitmap <= 16'b0000000000000000;
		15'h4ac3: char_row_bitmap <= 16'b0000000000000000;
		15'h4ac4: char_row_bitmap <= 16'b0011111100000000;
		15'h4ac5: char_row_bitmap <= 16'b0011111100000000;
		15'h4ac6: char_row_bitmap <= 16'b0011111100000000;
		15'h4ac7: char_row_bitmap <= 16'b0011111100000000;
		15'h4ac8: char_row_bitmap <= 16'b0000000000000000;
		15'h4ac9: char_row_bitmap <= 16'b0000000000000000;
		15'h4aca: char_row_bitmap <= 16'b0011111100111111;
		15'h4acb: char_row_bitmap <= 16'b0011111100111111;
		15'h4acc: char_row_bitmap <= 16'b0011111100111111;
		15'h4acd: char_row_bitmap <= 16'b0011111100111111;
		15'h4ace: char_row_bitmap <= 16'b0011111100111111;
		15'h4acf: char_row_bitmap <= 16'b0011111100111111;
		15'h4ad0: char_row_bitmap <= 16'b0000000000000000;
		15'h4ad1: char_row_bitmap <= 16'b0000000000000000;
		15'h4ad2: char_row_bitmap <= 16'b0011111100111111;
		15'h4ad3: char_row_bitmap <= 16'b0011111100111111;
		15'h4ad4: char_row_bitmap <= 16'b0011111100111111;
		15'h4ad5: char_row_bitmap <= 16'b0011111100111111;
		15'h4ad6: char_row_bitmap <= 16'b0000000000000000;
		15'h4ad7: char_row_bitmap <= 16'b0000000000000000;
		15'h4ad8: char_row_bitmap <= 16'b0000000000111111;
		15'h4ad9: char_row_bitmap <= 16'b0000000000111111;
		15'h4ada: char_row_bitmap <= 16'b0000000000111111;
		15'h4adb: char_row_bitmap <= 16'b0000000000111111;
		15'h4adc: char_row_bitmap <= 16'b0000000000000000;
		15'h4add: char_row_bitmap <= 16'b0000000000000000;
		15'h4ade: char_row_bitmap <= 16'b0011111100111111;
		15'h4adf: char_row_bitmap <= 16'b0011111100111111;
		15'h4ae0: char_row_bitmap <= 16'b0011111100111111;
		15'h4ae1: char_row_bitmap <= 16'b0011111100111111;
		15'h4ae2: char_row_bitmap <= 16'b0011111100111111;
		15'h4ae3: char_row_bitmap <= 16'b0011111100111111;
		15'h4ae4: char_row_bitmap <= 16'b0000000000000000;
		15'h4ae5: char_row_bitmap <= 16'b0000000000000000;
		15'h4ae6: char_row_bitmap <= 16'b0011111100111111;
		15'h4ae7: char_row_bitmap <= 16'b0011111100111111;
		15'h4ae8: char_row_bitmap <= 16'b0011111100111111;
		15'h4ae9: char_row_bitmap <= 16'b0011111100111111;
		15'h4aea: char_row_bitmap <= 16'b0000000000000000;
		15'h4aeb: char_row_bitmap <= 16'b0000000000000000;
		15'h4aec: char_row_bitmap <= 16'b0011111100111111;
		15'h4aed: char_row_bitmap <= 16'b0011111100111111;
		15'h4aee: char_row_bitmap <= 16'b0011111100111111;
		15'h4aef: char_row_bitmap <= 16'b0011111100111111;
		15'h4af0: char_row_bitmap <= 16'b0000000000000000;
		15'h4af1: char_row_bitmap <= 16'b0000000000000000;
		15'h4af2: char_row_bitmap <= 16'b0011111100111111;
		15'h4af3: char_row_bitmap <= 16'b0011111100111111;
		15'h4af4: char_row_bitmap <= 16'b0011111100111111;
		15'h4af5: char_row_bitmap <= 16'b0011111100111111;
		15'h4af6: char_row_bitmap <= 16'b0011111100111111;
		15'h4af7: char_row_bitmap <= 16'b0011111100111111;
		15'h4af8: char_row_bitmap <= 16'b0000000000000000;
		15'h4af9: char_row_bitmap <= 16'b0000000000000000;
		15'h4afa: char_row_bitmap <= 16'b0011111100111111;
		15'h4afb: char_row_bitmap <= 16'b0011111100111111;
		15'h4afc: char_row_bitmap <= 16'b0011111100111111;
		15'h4afd: char_row_bitmap <= 16'b0011111100111111;
		15'h4afe: char_row_bitmap <= 16'b0000000000000000;
		15'h4aff: char_row_bitmap <= 16'b0000000000000000;
		15'h4b00: char_row_bitmap <= 16'b0000000000000000;
		15'h4b01: char_row_bitmap <= 16'b0000000000000000;
		15'h4b02: char_row_bitmap <= 16'b0000000000000000;
		15'h4b03: char_row_bitmap <= 16'b0000000000000000;
		15'h4b04: char_row_bitmap <= 16'b0000000000000000;
		15'h4b05: char_row_bitmap <= 16'b0000000000000000;
		15'h4b06: char_row_bitmap <= 16'b0000000000000000;
		15'h4b07: char_row_bitmap <= 16'b0000000000000000;
		15'h4b08: char_row_bitmap <= 16'b0000000000000000;
		15'h4b09: char_row_bitmap <= 16'b0000000000000000;
		15'h4b0a: char_row_bitmap <= 16'b0000000000000000;
		15'h4b0b: char_row_bitmap <= 16'b0000000000000000;
		15'h4b0c: char_row_bitmap <= 16'b0000000000000000;
		15'h4b0d: char_row_bitmap <= 16'b0000000000000000;
		15'h4b0e: char_row_bitmap <= 16'b0000000000000000;
		15'h4b0f: char_row_bitmap <= 16'b0000000000000000;
		15'h4b10: char_row_bitmap <= 16'b0000000000000000;
		15'h4b11: char_row_bitmap <= 16'b0000000000000000;
		15'h4b12: char_row_bitmap <= 16'b0000000000000000;
		15'h4b13: char_row_bitmap <= 16'b0000000000000000;
		15'h4b14: char_row_bitmap <= 16'b1111111100000000;
		15'h4b15: char_row_bitmap <= 16'b1111111100000000;
		15'h4b16: char_row_bitmap <= 16'b1111111100000000;
		15'h4b17: char_row_bitmap <= 16'b1111111100000000;
		15'h4b18: char_row_bitmap <= 16'b1111111100000000;
		15'h4b19: char_row_bitmap <= 16'b1111111100000000;
		15'h4b1a: char_row_bitmap <= 16'b0000000000000000;
		15'h4b1b: char_row_bitmap <= 16'b0000000000000000;
		15'h4b1c: char_row_bitmap <= 16'b0000000000000000;
		15'h4b1d: char_row_bitmap <= 16'b0000000000000000;
		15'h4b1e: char_row_bitmap <= 16'b0000000000000000;
		15'h4b1f: char_row_bitmap <= 16'b0000000000000000;
		15'h4b20: char_row_bitmap <= 16'b0000000000000000;
		15'h4b21: char_row_bitmap <= 16'b0000000000000000;
		15'h4b22: char_row_bitmap <= 16'b0000000000000000;
		15'h4b23: char_row_bitmap <= 16'b0000000000000000;
		15'h4b24: char_row_bitmap <= 16'b0000000000000000;
		15'h4b25: char_row_bitmap <= 16'b0000000000000000;
		15'h4b26: char_row_bitmap <= 16'b0000000000000000;
		15'h4b27: char_row_bitmap <= 16'b0000000000000000;
		15'h4b28: char_row_bitmap <= 16'b0000000011111111;
		15'h4b29: char_row_bitmap <= 16'b0000000011111111;
		15'h4b2a: char_row_bitmap <= 16'b0000000011111111;
		15'h4b2b: char_row_bitmap <= 16'b0000000011111111;
		15'h4b2c: char_row_bitmap <= 16'b0000000011111111;
		15'h4b2d: char_row_bitmap <= 16'b0000000011111111;
		15'h4b2e: char_row_bitmap <= 16'b0000000000000000;
		15'h4b2f: char_row_bitmap <= 16'b0000000000000000;
		15'h4b30: char_row_bitmap <= 16'b0000000000000000;
		15'h4b31: char_row_bitmap <= 16'b0000000000000000;
		15'h4b32: char_row_bitmap <= 16'b0000000000000000;
		15'h4b33: char_row_bitmap <= 16'b0000000000000000;
		15'h4b34: char_row_bitmap <= 16'b0000000000000000;
		15'h4b35: char_row_bitmap <= 16'b0000000000000000;
		15'h4b36: char_row_bitmap <= 16'b0000000000000000;
		15'h4b37: char_row_bitmap <= 16'b0000000000000000;
		15'h4b38: char_row_bitmap <= 16'b0000000000000000;
		15'h4b39: char_row_bitmap <= 16'b0000000000000000;
		15'h4b3a: char_row_bitmap <= 16'b0000000000000000;
		15'h4b3b: char_row_bitmap <= 16'b0000000000000000;
		15'h4b3c: char_row_bitmap <= 16'b1111111111111111;
		15'h4b3d: char_row_bitmap <= 16'b1111111111111111;
		15'h4b3e: char_row_bitmap <= 16'b1111111111111111;
		15'h4b3f: char_row_bitmap <= 16'b1111111111111111;
		15'h4b40: char_row_bitmap <= 16'b1111111111111111;
		15'h4b41: char_row_bitmap <= 16'b1111111111111111;
		15'h4b42: char_row_bitmap <= 16'b0000000000000000;
		15'h4b43: char_row_bitmap <= 16'b0000000000000000;
		15'h4b44: char_row_bitmap <= 16'b0000000000000000;
		15'h4b45: char_row_bitmap <= 16'b0000000000000000;
		15'h4b46: char_row_bitmap <= 16'b0000000000000000;
		15'h4b47: char_row_bitmap <= 16'b0000000000000000;
		15'h4b48: char_row_bitmap <= 16'b0000000000000000;
		15'h4b49: char_row_bitmap <= 16'b0000000000000000;
		15'h4b4a: char_row_bitmap <= 16'b0000000000000000;
		15'h4b4b: char_row_bitmap <= 16'b0000000000000000;
		15'h4b4c: char_row_bitmap <= 16'b0000000000000000;
		15'h4b4d: char_row_bitmap <= 16'b0000000000000000;
		15'h4b4e: char_row_bitmap <= 16'b0000000000000000;
		15'h4b4f: char_row_bitmap <= 16'b0000000000000000;
		15'h4b50: char_row_bitmap <= 16'b0000000000000000;
		15'h4b51: char_row_bitmap <= 16'b0000000000000000;
		15'h4b52: char_row_bitmap <= 16'b0000000000000000;
		15'h4b53: char_row_bitmap <= 16'b0000000000000000;
		15'h4b54: char_row_bitmap <= 16'b0000000000000000;
		15'h4b55: char_row_bitmap <= 16'b0000000000000000;
		15'h4b56: char_row_bitmap <= 16'b1111111100000000;
		15'h4b57: char_row_bitmap <= 16'b1111111100000000;
		15'h4b58: char_row_bitmap <= 16'b1111111100000000;
		15'h4b59: char_row_bitmap <= 16'b1111111100000000;
		15'h4b5a: char_row_bitmap <= 16'b1111111100000000;
		15'h4b5b: char_row_bitmap <= 16'b1111111100000000;
		15'h4b5c: char_row_bitmap <= 16'b1111111100000000;
		15'h4b5d: char_row_bitmap <= 16'b1111111100000000;
		15'h4b5e: char_row_bitmap <= 16'b0000000000000000;
		15'h4b5f: char_row_bitmap <= 16'b0000000000000000;
		15'h4b60: char_row_bitmap <= 16'b0000000000000000;
		15'h4b61: char_row_bitmap <= 16'b0000000000000000;
		15'h4b62: char_row_bitmap <= 16'b0000000000000000;
		15'h4b63: char_row_bitmap <= 16'b0000000000000000;
		15'h4b64: char_row_bitmap <= 16'b1111111100000000;
		15'h4b65: char_row_bitmap <= 16'b1111111100000000;
		15'h4b66: char_row_bitmap <= 16'b1111111100000000;
		15'h4b67: char_row_bitmap <= 16'b1111111100000000;
		15'h4b68: char_row_bitmap <= 16'b1111111100000000;
		15'h4b69: char_row_bitmap <= 16'b1111111100000000;
		15'h4b6a: char_row_bitmap <= 16'b1111111100000000;
		15'h4b6b: char_row_bitmap <= 16'b1111111100000000;
		15'h4b6c: char_row_bitmap <= 16'b1111111100000000;
		15'h4b6d: char_row_bitmap <= 16'b1111111100000000;
		15'h4b6e: char_row_bitmap <= 16'b1111111100000000;
		15'h4b6f: char_row_bitmap <= 16'b1111111100000000;
		15'h4b70: char_row_bitmap <= 16'b1111111100000000;
		15'h4b71: char_row_bitmap <= 16'b1111111100000000;
		15'h4b72: char_row_bitmap <= 16'b0000000000000000;
		15'h4b73: char_row_bitmap <= 16'b0000000000000000;
		15'h4b74: char_row_bitmap <= 16'b0000000000000000;
		15'h4b75: char_row_bitmap <= 16'b0000000000000000;
		15'h4b76: char_row_bitmap <= 16'b0000000000000000;
		15'h4b77: char_row_bitmap <= 16'b0000000000000000;
		15'h4b78: char_row_bitmap <= 16'b0000000011111111;
		15'h4b79: char_row_bitmap <= 16'b0000000011111111;
		15'h4b7a: char_row_bitmap <= 16'b0000000011111111;
		15'h4b7b: char_row_bitmap <= 16'b0000000011111111;
		15'h4b7c: char_row_bitmap <= 16'b0000000011111111;
		15'h4b7d: char_row_bitmap <= 16'b0000000011111111;
		15'h4b7e: char_row_bitmap <= 16'b1111111100000000;
		15'h4b7f: char_row_bitmap <= 16'b1111111100000000;
		15'h4b80: char_row_bitmap <= 16'b1111111100000000;
		15'h4b81: char_row_bitmap <= 16'b1111111100000000;
		15'h4b82: char_row_bitmap <= 16'b1111111100000000;
		15'h4b83: char_row_bitmap <= 16'b1111111100000000;
		15'h4b84: char_row_bitmap <= 16'b1111111100000000;
		15'h4b85: char_row_bitmap <= 16'b1111111100000000;
		15'h4b86: char_row_bitmap <= 16'b0000000000000000;
		15'h4b87: char_row_bitmap <= 16'b0000000000000000;
		15'h4b88: char_row_bitmap <= 16'b0000000000000000;
		15'h4b89: char_row_bitmap <= 16'b0000000000000000;
		15'h4b8a: char_row_bitmap <= 16'b0000000000000000;
		15'h4b8b: char_row_bitmap <= 16'b0000000000000000;
		15'h4b8c: char_row_bitmap <= 16'b1111111111111111;
		15'h4b8d: char_row_bitmap <= 16'b1111111111111111;
		15'h4b8e: char_row_bitmap <= 16'b1111111111111111;
		15'h4b8f: char_row_bitmap <= 16'b1111111111111111;
		15'h4b90: char_row_bitmap <= 16'b1111111111111111;
		15'h4b91: char_row_bitmap <= 16'b1111111111111111;
		15'h4b92: char_row_bitmap <= 16'b1111111100000000;
		15'h4b93: char_row_bitmap <= 16'b1111111100000000;
		15'h4b94: char_row_bitmap <= 16'b1111111100000000;
		15'h4b95: char_row_bitmap <= 16'b1111111100000000;
		15'h4b96: char_row_bitmap <= 16'b1111111100000000;
		15'h4b97: char_row_bitmap <= 16'b1111111100000000;
		15'h4b98: char_row_bitmap <= 16'b1111111100000000;
		15'h4b99: char_row_bitmap <= 16'b1111111100000000;
		15'h4b9a: char_row_bitmap <= 16'b0000000000000000;
		15'h4b9b: char_row_bitmap <= 16'b0000000000000000;
		15'h4b9c: char_row_bitmap <= 16'b0000000000000000;
		15'h4b9d: char_row_bitmap <= 16'b0000000000000000;
		15'h4b9e: char_row_bitmap <= 16'b0000000000000000;
		15'h4b9f: char_row_bitmap <= 16'b0000000000000000;
		15'h4ba0: char_row_bitmap <= 16'b0000000000000000;
		15'h4ba1: char_row_bitmap <= 16'b0000000000000000;
		15'h4ba2: char_row_bitmap <= 16'b0000000000000000;
		15'h4ba3: char_row_bitmap <= 16'b0000000000000000;
		15'h4ba4: char_row_bitmap <= 16'b0000000000000000;
		15'h4ba5: char_row_bitmap <= 16'b0000000000000000;
		15'h4ba6: char_row_bitmap <= 16'b0000000011111111;
		15'h4ba7: char_row_bitmap <= 16'b0000000011111111;
		15'h4ba8: char_row_bitmap <= 16'b0000000011111111;
		15'h4ba9: char_row_bitmap <= 16'b0000000011111111;
		15'h4baa: char_row_bitmap <= 16'b0000000011111111;
		15'h4bab: char_row_bitmap <= 16'b0000000011111111;
		15'h4bac: char_row_bitmap <= 16'b0000000011111111;
		15'h4bad: char_row_bitmap <= 16'b0000000011111111;
		15'h4bae: char_row_bitmap <= 16'b0000000000000000;
		15'h4baf: char_row_bitmap <= 16'b0000000000000000;
		15'h4bb0: char_row_bitmap <= 16'b0000000000000000;
		15'h4bb1: char_row_bitmap <= 16'b0000000000000000;
		15'h4bb2: char_row_bitmap <= 16'b0000000000000000;
		15'h4bb3: char_row_bitmap <= 16'b0000000000000000;
		15'h4bb4: char_row_bitmap <= 16'b1111111100000000;
		15'h4bb5: char_row_bitmap <= 16'b1111111100000000;
		15'h4bb6: char_row_bitmap <= 16'b1111111100000000;
		15'h4bb7: char_row_bitmap <= 16'b1111111100000000;
		15'h4bb8: char_row_bitmap <= 16'b1111111100000000;
		15'h4bb9: char_row_bitmap <= 16'b1111111100000000;
		15'h4bba: char_row_bitmap <= 16'b0000000011111111;
		15'h4bbb: char_row_bitmap <= 16'b0000000011111111;
		15'h4bbc: char_row_bitmap <= 16'b0000000011111111;
		15'h4bbd: char_row_bitmap <= 16'b0000000011111111;
		15'h4bbe: char_row_bitmap <= 16'b0000000011111111;
		15'h4bbf: char_row_bitmap <= 16'b0000000011111111;
		15'h4bc0: char_row_bitmap <= 16'b0000000011111111;
		15'h4bc1: char_row_bitmap <= 16'b0000000011111111;
		15'h4bc2: char_row_bitmap <= 16'b0000000000000000;
		15'h4bc3: char_row_bitmap <= 16'b0000000000000000;
		15'h4bc4: char_row_bitmap <= 16'b0000000000000000;
		15'h4bc5: char_row_bitmap <= 16'b0000000000000000;
		15'h4bc6: char_row_bitmap <= 16'b0000000000000000;
		15'h4bc7: char_row_bitmap <= 16'b0000000000000000;
		15'h4bc8: char_row_bitmap <= 16'b0000000011111111;
		15'h4bc9: char_row_bitmap <= 16'b0000000011111111;
		15'h4bca: char_row_bitmap <= 16'b0000000011111111;
		15'h4bcb: char_row_bitmap <= 16'b0000000011111111;
		15'h4bcc: char_row_bitmap <= 16'b0000000011111111;
		15'h4bcd: char_row_bitmap <= 16'b0000000011111111;
		15'h4bce: char_row_bitmap <= 16'b0000000011111111;
		15'h4bcf: char_row_bitmap <= 16'b0000000011111111;
		15'h4bd0: char_row_bitmap <= 16'b0000000011111111;
		15'h4bd1: char_row_bitmap <= 16'b0000000011111111;
		15'h4bd2: char_row_bitmap <= 16'b0000000011111111;
		15'h4bd3: char_row_bitmap <= 16'b0000000011111111;
		15'h4bd4: char_row_bitmap <= 16'b0000000011111111;
		15'h4bd5: char_row_bitmap <= 16'b0000000011111111;
		15'h4bd6: char_row_bitmap <= 16'b0000000000000000;
		15'h4bd7: char_row_bitmap <= 16'b0000000000000000;
		15'h4bd8: char_row_bitmap <= 16'b0000000000000000;
		15'h4bd9: char_row_bitmap <= 16'b0000000000000000;
		15'h4bda: char_row_bitmap <= 16'b0000000000000000;
		15'h4bdb: char_row_bitmap <= 16'b0000000000000000;
		15'h4bdc: char_row_bitmap <= 16'b1111111111111111;
		15'h4bdd: char_row_bitmap <= 16'b1111111111111111;
		15'h4bde: char_row_bitmap <= 16'b1111111111111111;
		15'h4bdf: char_row_bitmap <= 16'b1111111111111111;
		15'h4be0: char_row_bitmap <= 16'b1111111111111111;
		15'h4be1: char_row_bitmap <= 16'b1111111111111111;
		15'h4be2: char_row_bitmap <= 16'b0000000011111111;
		15'h4be3: char_row_bitmap <= 16'b0000000011111111;
		15'h4be4: char_row_bitmap <= 16'b0000000011111111;
		15'h4be5: char_row_bitmap <= 16'b0000000011111111;
		15'h4be6: char_row_bitmap <= 16'b0000000011111111;
		15'h4be7: char_row_bitmap <= 16'b0000000011111111;
		15'h4be8: char_row_bitmap <= 16'b0000000011111111;
		15'h4be9: char_row_bitmap <= 16'b0000000011111111;
		15'h4bea: char_row_bitmap <= 16'b0000000000000000;
		15'h4beb: char_row_bitmap <= 16'b0000000000000000;
		15'h4bec: char_row_bitmap <= 16'b0000000000000000;
		15'h4bed: char_row_bitmap <= 16'b0000000000000000;
		15'h4bee: char_row_bitmap <= 16'b0000000000000000;
		15'h4bef: char_row_bitmap <= 16'b0000000000000000;
		15'h4bf0: char_row_bitmap <= 16'b0000000000000000;
		15'h4bf1: char_row_bitmap <= 16'b0000000000000000;
		15'h4bf2: char_row_bitmap <= 16'b0000000000000000;
		15'h4bf3: char_row_bitmap <= 16'b0000000000000000;
		15'h4bf4: char_row_bitmap <= 16'b0000000000000000;
		15'h4bf5: char_row_bitmap <= 16'b0000000000000000;
		15'h4bf6: char_row_bitmap <= 16'b1111111111111111;
		15'h4bf7: char_row_bitmap <= 16'b1111111111111111;
		15'h4bf8: char_row_bitmap <= 16'b1111111111111111;
		15'h4bf9: char_row_bitmap <= 16'b1111111111111111;
		15'h4bfa: char_row_bitmap <= 16'b1111111111111111;
		15'h4bfb: char_row_bitmap <= 16'b1111111111111111;
		15'h4bfc: char_row_bitmap <= 16'b1111111111111111;
		15'h4bfd: char_row_bitmap <= 16'b1111111111111111;
		15'h4bfe: char_row_bitmap <= 16'b0000000000000000;
		15'h4bff: char_row_bitmap <= 16'b0000000000000000;
		15'h4c00: char_row_bitmap <= 16'b0000000000000000;
		15'h4c01: char_row_bitmap <= 16'b0000000000000000;
		15'h4c02: char_row_bitmap <= 16'b0000000000000000;
		15'h4c03: char_row_bitmap <= 16'b0000000000000000;
		15'h4c04: char_row_bitmap <= 16'b1111111100000000;
		15'h4c05: char_row_bitmap <= 16'b1111111100000000;
		15'h4c06: char_row_bitmap <= 16'b1111111100000000;
		15'h4c07: char_row_bitmap <= 16'b1111111100000000;
		15'h4c08: char_row_bitmap <= 16'b1111111100000000;
		15'h4c09: char_row_bitmap <= 16'b1111111100000000;
		15'h4c0a: char_row_bitmap <= 16'b1111111111111111;
		15'h4c0b: char_row_bitmap <= 16'b1111111111111111;
		15'h4c0c: char_row_bitmap <= 16'b1111111111111111;
		15'h4c0d: char_row_bitmap <= 16'b1111111111111111;
		15'h4c0e: char_row_bitmap <= 16'b1111111111111111;
		15'h4c0f: char_row_bitmap <= 16'b1111111111111111;
		15'h4c10: char_row_bitmap <= 16'b1111111111111111;
		15'h4c11: char_row_bitmap <= 16'b1111111111111111;
		15'h4c12: char_row_bitmap <= 16'b0000000000000000;
		15'h4c13: char_row_bitmap <= 16'b0000000000000000;
		15'h4c14: char_row_bitmap <= 16'b0000000000000000;
		15'h4c15: char_row_bitmap <= 16'b0000000000000000;
		15'h4c16: char_row_bitmap <= 16'b0000000000000000;
		15'h4c17: char_row_bitmap <= 16'b0000000000000000;
		15'h4c18: char_row_bitmap <= 16'b0000000011111111;
		15'h4c19: char_row_bitmap <= 16'b0000000011111111;
		15'h4c1a: char_row_bitmap <= 16'b0000000011111111;
		15'h4c1b: char_row_bitmap <= 16'b0000000011111111;
		15'h4c1c: char_row_bitmap <= 16'b0000000011111111;
		15'h4c1d: char_row_bitmap <= 16'b0000000011111111;
		15'h4c1e: char_row_bitmap <= 16'b1111111111111111;
		15'h4c1f: char_row_bitmap <= 16'b1111111111111111;
		15'h4c20: char_row_bitmap <= 16'b1111111111111111;
		15'h4c21: char_row_bitmap <= 16'b1111111111111111;
		15'h4c22: char_row_bitmap <= 16'b1111111111111111;
		15'h4c23: char_row_bitmap <= 16'b1111111111111111;
		15'h4c24: char_row_bitmap <= 16'b1111111111111111;
		15'h4c25: char_row_bitmap <= 16'b1111111111111111;
		15'h4c26: char_row_bitmap <= 16'b0000000000000000;
		15'h4c27: char_row_bitmap <= 16'b0000000000000000;
		15'h4c28: char_row_bitmap <= 16'b0000000000000000;
		15'h4c29: char_row_bitmap <= 16'b0000000000000000;
		15'h4c2a: char_row_bitmap <= 16'b0000000000000000;
		15'h4c2b: char_row_bitmap <= 16'b0000000000000000;
		15'h4c2c: char_row_bitmap <= 16'b1111111111111111;
		15'h4c2d: char_row_bitmap <= 16'b1111111111111111;
		15'h4c2e: char_row_bitmap <= 16'b1111111111111111;
		15'h4c2f: char_row_bitmap <= 16'b1111111111111111;
		15'h4c30: char_row_bitmap <= 16'b1111111111111111;
		15'h4c31: char_row_bitmap <= 16'b1111111111111111;
		15'h4c32: char_row_bitmap <= 16'b1111111111111111;
		15'h4c33: char_row_bitmap <= 16'b1111111111111111;
		15'h4c34: char_row_bitmap <= 16'b1111111111111111;
		15'h4c35: char_row_bitmap <= 16'b1111111111111111;
		15'h4c36: char_row_bitmap <= 16'b1111111111111111;
		15'h4c37: char_row_bitmap <= 16'b1111111111111111;
		15'h4c38: char_row_bitmap <= 16'b1111111111111111;
		15'h4c39: char_row_bitmap <= 16'b1111111111111111;
		15'h4c3a: char_row_bitmap <= 16'b0000000000000000;
		15'h4c3b: char_row_bitmap <= 16'b0000000000000000;
		15'h4c3c: char_row_bitmap <= 16'b0000000000000000;
		15'h4c3d: char_row_bitmap <= 16'b0000000000000000;
		15'h4c3e: char_row_bitmap <= 16'b0000000000000000;
		15'h4c3f: char_row_bitmap <= 16'b0000000000000000;
		15'h4c40: char_row_bitmap <= 16'b0000000000000000;
		15'h4c41: char_row_bitmap <= 16'b0000000000000000;
		15'h4c42: char_row_bitmap <= 16'b0000000000000000;
		15'h4c43: char_row_bitmap <= 16'b0000000000000000;
		15'h4c44: char_row_bitmap <= 16'b0000000000000000;
		15'h4c45: char_row_bitmap <= 16'b0000000000000000;
		15'h4c46: char_row_bitmap <= 16'b0000000000000000;
		15'h4c47: char_row_bitmap <= 16'b0000000000000000;
		15'h4c48: char_row_bitmap <= 16'b0000000000000000;
		15'h4c49: char_row_bitmap <= 16'b0000000000000000;
		15'h4c4a: char_row_bitmap <= 16'b0000000000000000;
		15'h4c4b: char_row_bitmap <= 16'b0000000000000000;
		15'h4c4c: char_row_bitmap <= 16'b0000000000000000;
		15'h4c4d: char_row_bitmap <= 16'b0000000000000000;
		15'h4c4e: char_row_bitmap <= 16'b1111111100000000;
		15'h4c4f: char_row_bitmap <= 16'b1111111100000000;
		15'h4c50: char_row_bitmap <= 16'b1111111100000000;
		15'h4c51: char_row_bitmap <= 16'b1111111100000000;
		15'h4c52: char_row_bitmap <= 16'b1111111100000000;
		15'h4c53: char_row_bitmap <= 16'b1111111100000000;
		15'h4c54: char_row_bitmap <= 16'b1111111100000000;
		15'h4c55: char_row_bitmap <= 16'b1111111100000000;
		15'h4c56: char_row_bitmap <= 16'b1111111100000000;
		15'h4c57: char_row_bitmap <= 16'b1111111100000000;
		15'h4c58: char_row_bitmap <= 16'b1111111100000000;
		15'h4c59: char_row_bitmap <= 16'b1111111100000000;
		15'h4c5a: char_row_bitmap <= 16'b0000000000000000;
		15'h4c5b: char_row_bitmap <= 16'b0000000000000000;
		15'h4c5c: char_row_bitmap <= 16'b0000000000000000;
		15'h4c5d: char_row_bitmap <= 16'b0000000000000000;
		15'h4c5e: char_row_bitmap <= 16'b0000000000000000;
		15'h4c5f: char_row_bitmap <= 16'b0000000000000000;
		15'h4c60: char_row_bitmap <= 16'b0000000000000000;
		15'h4c61: char_row_bitmap <= 16'b0000000000000000;
		15'h4c62: char_row_bitmap <= 16'b1111111100000000;
		15'h4c63: char_row_bitmap <= 16'b1111111100000000;
		15'h4c64: char_row_bitmap <= 16'b1111111100000000;
		15'h4c65: char_row_bitmap <= 16'b1111111100000000;
		15'h4c66: char_row_bitmap <= 16'b1111111100000000;
		15'h4c67: char_row_bitmap <= 16'b1111111100000000;
		15'h4c68: char_row_bitmap <= 16'b0000000011111111;
		15'h4c69: char_row_bitmap <= 16'b0000000011111111;
		15'h4c6a: char_row_bitmap <= 16'b0000000011111111;
		15'h4c6b: char_row_bitmap <= 16'b0000000011111111;
		15'h4c6c: char_row_bitmap <= 16'b0000000011111111;
		15'h4c6d: char_row_bitmap <= 16'b0000000011111111;
		15'h4c6e: char_row_bitmap <= 16'b0000000000000000;
		15'h4c6f: char_row_bitmap <= 16'b0000000000000000;
		15'h4c70: char_row_bitmap <= 16'b0000000000000000;
		15'h4c71: char_row_bitmap <= 16'b0000000000000000;
		15'h4c72: char_row_bitmap <= 16'b0000000000000000;
		15'h4c73: char_row_bitmap <= 16'b0000000000000000;
		15'h4c74: char_row_bitmap <= 16'b0000000000000000;
		15'h4c75: char_row_bitmap <= 16'b0000000000000000;
		15'h4c76: char_row_bitmap <= 16'b1111111100000000;
		15'h4c77: char_row_bitmap <= 16'b1111111100000000;
		15'h4c78: char_row_bitmap <= 16'b1111111100000000;
		15'h4c79: char_row_bitmap <= 16'b1111111100000000;
		15'h4c7a: char_row_bitmap <= 16'b1111111100000000;
		15'h4c7b: char_row_bitmap <= 16'b1111111100000000;
		15'h4c7c: char_row_bitmap <= 16'b1111111111111111;
		15'h4c7d: char_row_bitmap <= 16'b1111111111111111;
		15'h4c7e: char_row_bitmap <= 16'b1111111111111111;
		15'h4c7f: char_row_bitmap <= 16'b1111111111111111;
		15'h4c80: char_row_bitmap <= 16'b1111111111111111;
		15'h4c81: char_row_bitmap <= 16'b1111111111111111;
		15'h4c82: char_row_bitmap <= 16'b0000000000000000;
		15'h4c83: char_row_bitmap <= 16'b0000000000000000;
		15'h4c84: char_row_bitmap <= 16'b0000000000000000;
		15'h4c85: char_row_bitmap <= 16'b0000000000000000;
		15'h4c86: char_row_bitmap <= 16'b0000000000000000;
		15'h4c87: char_row_bitmap <= 16'b0000000000000000;
		15'h4c88: char_row_bitmap <= 16'b0000000000000000;
		15'h4c89: char_row_bitmap <= 16'b0000000000000000;
		15'h4c8a: char_row_bitmap <= 16'b1111111100000000;
		15'h4c8b: char_row_bitmap <= 16'b1111111100000000;
		15'h4c8c: char_row_bitmap <= 16'b1111111100000000;
		15'h4c8d: char_row_bitmap <= 16'b1111111100000000;
		15'h4c8e: char_row_bitmap <= 16'b1111111100000000;
		15'h4c8f: char_row_bitmap <= 16'b1111111100000000;
		15'h4c90: char_row_bitmap <= 16'b0000000000000000;
		15'h4c91: char_row_bitmap <= 16'b0000000000000000;
		15'h4c92: char_row_bitmap <= 16'b0000000000000000;
		15'h4c93: char_row_bitmap <= 16'b0000000000000000;
		15'h4c94: char_row_bitmap <= 16'b0000000000000000;
		15'h4c95: char_row_bitmap <= 16'b0000000000000000;
		15'h4c96: char_row_bitmap <= 16'b1111111100000000;
		15'h4c97: char_row_bitmap <= 16'b1111111100000000;
		15'h4c98: char_row_bitmap <= 16'b1111111100000000;
		15'h4c99: char_row_bitmap <= 16'b1111111100000000;
		15'h4c9a: char_row_bitmap <= 16'b1111111100000000;
		15'h4c9b: char_row_bitmap <= 16'b1111111100000000;
		15'h4c9c: char_row_bitmap <= 16'b1111111100000000;
		15'h4c9d: char_row_bitmap <= 16'b1111111100000000;
		15'h4c9e: char_row_bitmap <= 16'b1111111100000000;
		15'h4c9f: char_row_bitmap <= 16'b1111111100000000;
		15'h4ca0: char_row_bitmap <= 16'b1111111100000000;
		15'h4ca1: char_row_bitmap <= 16'b1111111100000000;
		15'h4ca2: char_row_bitmap <= 16'b1111111100000000;
		15'h4ca3: char_row_bitmap <= 16'b1111111100000000;
		15'h4ca4: char_row_bitmap <= 16'b1111111100000000;
		15'h4ca5: char_row_bitmap <= 16'b1111111100000000;
		15'h4ca6: char_row_bitmap <= 16'b1111111100000000;
		15'h4ca7: char_row_bitmap <= 16'b1111111100000000;
		15'h4ca8: char_row_bitmap <= 16'b1111111100000000;
		15'h4ca9: char_row_bitmap <= 16'b1111111100000000;
		15'h4caa: char_row_bitmap <= 16'b1111111100000000;
		15'h4cab: char_row_bitmap <= 16'b1111111100000000;
		15'h4cac: char_row_bitmap <= 16'b1111111100000000;
		15'h4cad: char_row_bitmap <= 16'b1111111100000000;
		15'h4cae: char_row_bitmap <= 16'b1111111100000000;
		15'h4caf: char_row_bitmap <= 16'b1111111100000000;
		15'h4cb0: char_row_bitmap <= 16'b1111111100000000;
		15'h4cb1: char_row_bitmap <= 16'b1111111100000000;
		15'h4cb2: char_row_bitmap <= 16'b1111111100000000;
		15'h4cb3: char_row_bitmap <= 16'b1111111100000000;
		15'h4cb4: char_row_bitmap <= 16'b1111111100000000;
		15'h4cb5: char_row_bitmap <= 16'b1111111100000000;
		15'h4cb6: char_row_bitmap <= 16'b1111111100000000;
		15'h4cb7: char_row_bitmap <= 16'b1111111100000000;
		15'h4cb8: char_row_bitmap <= 16'b0000000011111111;
		15'h4cb9: char_row_bitmap <= 16'b0000000011111111;
		15'h4cba: char_row_bitmap <= 16'b0000000011111111;
		15'h4cbb: char_row_bitmap <= 16'b0000000011111111;
		15'h4cbc: char_row_bitmap <= 16'b0000000011111111;
		15'h4cbd: char_row_bitmap <= 16'b0000000011111111;
		15'h4cbe: char_row_bitmap <= 16'b1111111100000000;
		15'h4cbf: char_row_bitmap <= 16'b1111111100000000;
		15'h4cc0: char_row_bitmap <= 16'b1111111100000000;
		15'h4cc1: char_row_bitmap <= 16'b1111111100000000;
		15'h4cc2: char_row_bitmap <= 16'b1111111100000000;
		15'h4cc3: char_row_bitmap <= 16'b1111111100000000;
		15'h4cc4: char_row_bitmap <= 16'b1111111100000000;
		15'h4cc5: char_row_bitmap <= 16'b1111111100000000;
		15'h4cc6: char_row_bitmap <= 16'b1111111100000000;
		15'h4cc7: char_row_bitmap <= 16'b1111111100000000;
		15'h4cc8: char_row_bitmap <= 16'b1111111100000000;
		15'h4cc9: char_row_bitmap <= 16'b1111111100000000;
		15'h4cca: char_row_bitmap <= 16'b1111111100000000;
		15'h4ccb: char_row_bitmap <= 16'b1111111100000000;
		15'h4ccc: char_row_bitmap <= 16'b1111111111111111;
		15'h4ccd: char_row_bitmap <= 16'b1111111111111111;
		15'h4cce: char_row_bitmap <= 16'b1111111111111111;
		15'h4ccf: char_row_bitmap <= 16'b1111111111111111;
		15'h4cd0: char_row_bitmap <= 16'b1111111111111111;
		15'h4cd1: char_row_bitmap <= 16'b1111111111111111;
		15'h4cd2: char_row_bitmap <= 16'b1111111100000000;
		15'h4cd3: char_row_bitmap <= 16'b1111111100000000;
		15'h4cd4: char_row_bitmap <= 16'b1111111100000000;
		15'h4cd5: char_row_bitmap <= 16'b1111111100000000;
		15'h4cd6: char_row_bitmap <= 16'b1111111100000000;
		15'h4cd7: char_row_bitmap <= 16'b1111111100000000;
		15'h4cd8: char_row_bitmap <= 16'b1111111100000000;
		15'h4cd9: char_row_bitmap <= 16'b1111111100000000;
		15'h4cda: char_row_bitmap <= 16'b1111111100000000;
		15'h4cdb: char_row_bitmap <= 16'b1111111100000000;
		15'h4cdc: char_row_bitmap <= 16'b1111111100000000;
		15'h4cdd: char_row_bitmap <= 16'b1111111100000000;
		15'h4cde: char_row_bitmap <= 16'b1111111100000000;
		15'h4cdf: char_row_bitmap <= 16'b1111111100000000;
		15'h4ce0: char_row_bitmap <= 16'b0000000000000000;
		15'h4ce1: char_row_bitmap <= 16'b0000000000000000;
		15'h4ce2: char_row_bitmap <= 16'b0000000000000000;
		15'h4ce3: char_row_bitmap <= 16'b0000000000000000;
		15'h4ce4: char_row_bitmap <= 16'b0000000000000000;
		15'h4ce5: char_row_bitmap <= 16'b0000000000000000;
		15'h4ce6: char_row_bitmap <= 16'b0000000011111111;
		15'h4ce7: char_row_bitmap <= 16'b0000000011111111;
		15'h4ce8: char_row_bitmap <= 16'b0000000011111111;
		15'h4ce9: char_row_bitmap <= 16'b0000000011111111;
		15'h4cea: char_row_bitmap <= 16'b0000000011111111;
		15'h4ceb: char_row_bitmap <= 16'b0000000011111111;
		15'h4cec: char_row_bitmap <= 16'b0000000011111111;
		15'h4ced: char_row_bitmap <= 16'b0000000011111111;
		15'h4cee: char_row_bitmap <= 16'b1111111100000000;
		15'h4cef: char_row_bitmap <= 16'b1111111100000000;
		15'h4cf0: char_row_bitmap <= 16'b1111111100000000;
		15'h4cf1: char_row_bitmap <= 16'b1111111100000000;
		15'h4cf2: char_row_bitmap <= 16'b1111111100000000;
		15'h4cf3: char_row_bitmap <= 16'b1111111100000000;
		15'h4cf4: char_row_bitmap <= 16'b1111111100000000;
		15'h4cf5: char_row_bitmap <= 16'b1111111100000000;
		15'h4cf6: char_row_bitmap <= 16'b1111111100000000;
		15'h4cf7: char_row_bitmap <= 16'b1111111100000000;
		15'h4cf8: char_row_bitmap <= 16'b1111111100000000;
		15'h4cf9: char_row_bitmap <= 16'b1111111100000000;
		15'h4cfa: char_row_bitmap <= 16'b0000000011111111;
		15'h4cfb: char_row_bitmap <= 16'b0000000011111111;
		15'h4cfc: char_row_bitmap <= 16'b0000000011111111;
		15'h4cfd: char_row_bitmap <= 16'b0000000011111111;
		15'h4cfe: char_row_bitmap <= 16'b0000000011111111;
		15'h4cff: char_row_bitmap <= 16'b0000000011111111;
		15'h4d00: char_row_bitmap <= 16'b0000000011111111;
		15'h4d01: char_row_bitmap <= 16'b0000000011111111;
		15'h4d02: char_row_bitmap <= 16'b1111111100000000;
		15'h4d03: char_row_bitmap <= 16'b1111111100000000;
		15'h4d04: char_row_bitmap <= 16'b1111111100000000;
		15'h4d05: char_row_bitmap <= 16'b1111111100000000;
		15'h4d06: char_row_bitmap <= 16'b1111111100000000;
		15'h4d07: char_row_bitmap <= 16'b1111111100000000;
		15'h4d08: char_row_bitmap <= 16'b0000000011111111;
		15'h4d09: char_row_bitmap <= 16'b0000000011111111;
		15'h4d0a: char_row_bitmap <= 16'b0000000011111111;
		15'h4d0b: char_row_bitmap <= 16'b0000000011111111;
		15'h4d0c: char_row_bitmap <= 16'b0000000011111111;
		15'h4d0d: char_row_bitmap <= 16'b0000000011111111;
		15'h4d0e: char_row_bitmap <= 16'b0000000011111111;
		15'h4d0f: char_row_bitmap <= 16'b0000000011111111;
		15'h4d10: char_row_bitmap <= 16'b0000000011111111;
		15'h4d11: char_row_bitmap <= 16'b0000000011111111;
		15'h4d12: char_row_bitmap <= 16'b0000000011111111;
		15'h4d13: char_row_bitmap <= 16'b0000000011111111;
		15'h4d14: char_row_bitmap <= 16'b0000000011111111;
		15'h4d15: char_row_bitmap <= 16'b0000000011111111;
		15'h4d16: char_row_bitmap <= 16'b1111111100000000;
		15'h4d17: char_row_bitmap <= 16'b1111111100000000;
		15'h4d18: char_row_bitmap <= 16'b1111111100000000;
		15'h4d19: char_row_bitmap <= 16'b1111111100000000;
		15'h4d1a: char_row_bitmap <= 16'b1111111100000000;
		15'h4d1b: char_row_bitmap <= 16'b1111111100000000;
		15'h4d1c: char_row_bitmap <= 16'b1111111111111111;
		15'h4d1d: char_row_bitmap <= 16'b1111111111111111;
		15'h4d1e: char_row_bitmap <= 16'b1111111111111111;
		15'h4d1f: char_row_bitmap <= 16'b1111111111111111;
		15'h4d20: char_row_bitmap <= 16'b1111111111111111;
		15'h4d21: char_row_bitmap <= 16'b1111111111111111;
		15'h4d22: char_row_bitmap <= 16'b0000000011111111;
		15'h4d23: char_row_bitmap <= 16'b0000000011111111;
		15'h4d24: char_row_bitmap <= 16'b0000000011111111;
		15'h4d25: char_row_bitmap <= 16'b0000000011111111;
		15'h4d26: char_row_bitmap <= 16'b0000000011111111;
		15'h4d27: char_row_bitmap <= 16'b0000000011111111;
		15'h4d28: char_row_bitmap <= 16'b0000000011111111;
		15'h4d29: char_row_bitmap <= 16'b0000000011111111;
		15'h4d2a: char_row_bitmap <= 16'b1111111100000000;
		15'h4d2b: char_row_bitmap <= 16'b1111111100000000;
		15'h4d2c: char_row_bitmap <= 16'b1111111100000000;
		15'h4d2d: char_row_bitmap <= 16'b1111111100000000;
		15'h4d2e: char_row_bitmap <= 16'b1111111100000000;
		15'h4d2f: char_row_bitmap <= 16'b1111111100000000;
		15'h4d30: char_row_bitmap <= 16'b0000000000000000;
		15'h4d31: char_row_bitmap <= 16'b0000000000000000;
		15'h4d32: char_row_bitmap <= 16'b0000000000000000;
		15'h4d33: char_row_bitmap <= 16'b0000000000000000;
		15'h4d34: char_row_bitmap <= 16'b0000000000000000;
		15'h4d35: char_row_bitmap <= 16'b0000000000000000;
		15'h4d36: char_row_bitmap <= 16'b1111111111111111;
		15'h4d37: char_row_bitmap <= 16'b1111111111111111;
		15'h4d38: char_row_bitmap <= 16'b1111111111111111;
		15'h4d39: char_row_bitmap <= 16'b1111111111111111;
		15'h4d3a: char_row_bitmap <= 16'b1111111111111111;
		15'h4d3b: char_row_bitmap <= 16'b1111111111111111;
		15'h4d3c: char_row_bitmap <= 16'b1111111111111111;
		15'h4d3d: char_row_bitmap <= 16'b1111111111111111;
		15'h4d3e: char_row_bitmap <= 16'b1111111100000000;
		15'h4d3f: char_row_bitmap <= 16'b1111111100000000;
		15'h4d40: char_row_bitmap <= 16'b1111111100000000;
		15'h4d41: char_row_bitmap <= 16'b1111111100000000;
		15'h4d42: char_row_bitmap <= 16'b1111111100000000;
		15'h4d43: char_row_bitmap <= 16'b1111111100000000;
		15'h4d44: char_row_bitmap <= 16'b1111111100000000;
		15'h4d45: char_row_bitmap <= 16'b1111111100000000;
		15'h4d46: char_row_bitmap <= 16'b1111111100000000;
		15'h4d47: char_row_bitmap <= 16'b1111111100000000;
		15'h4d48: char_row_bitmap <= 16'b1111111100000000;
		15'h4d49: char_row_bitmap <= 16'b1111111100000000;
		15'h4d4a: char_row_bitmap <= 16'b1111111111111111;
		15'h4d4b: char_row_bitmap <= 16'b1111111111111111;
		15'h4d4c: char_row_bitmap <= 16'b1111111111111111;
		15'h4d4d: char_row_bitmap <= 16'b1111111111111111;
		15'h4d4e: char_row_bitmap <= 16'b1111111111111111;
		15'h4d4f: char_row_bitmap <= 16'b1111111111111111;
		15'h4d50: char_row_bitmap <= 16'b1111111111111111;
		15'h4d51: char_row_bitmap <= 16'b1111111111111111;
		15'h4d52: char_row_bitmap <= 16'b1111111100000000;
		15'h4d53: char_row_bitmap <= 16'b1111111100000000;
		15'h4d54: char_row_bitmap <= 16'b1111111100000000;
		15'h4d55: char_row_bitmap <= 16'b1111111100000000;
		15'h4d56: char_row_bitmap <= 16'b1111111100000000;
		15'h4d57: char_row_bitmap <= 16'b1111111100000000;
		15'h4d58: char_row_bitmap <= 16'b0000000011111111;
		15'h4d59: char_row_bitmap <= 16'b0000000011111111;
		15'h4d5a: char_row_bitmap <= 16'b0000000011111111;
		15'h4d5b: char_row_bitmap <= 16'b0000000011111111;
		15'h4d5c: char_row_bitmap <= 16'b0000000011111111;
		15'h4d5d: char_row_bitmap <= 16'b0000000011111111;
		15'h4d5e: char_row_bitmap <= 16'b1111111111111111;
		15'h4d5f: char_row_bitmap <= 16'b1111111111111111;
		15'h4d60: char_row_bitmap <= 16'b1111111111111111;
		15'h4d61: char_row_bitmap <= 16'b1111111111111111;
		15'h4d62: char_row_bitmap <= 16'b1111111111111111;
		15'h4d63: char_row_bitmap <= 16'b1111111111111111;
		15'h4d64: char_row_bitmap <= 16'b1111111111111111;
		15'h4d65: char_row_bitmap <= 16'b1111111111111111;
		15'h4d66: char_row_bitmap <= 16'b1111111100000000;
		15'h4d67: char_row_bitmap <= 16'b1111111100000000;
		15'h4d68: char_row_bitmap <= 16'b1111111100000000;
		15'h4d69: char_row_bitmap <= 16'b1111111100000000;
		15'h4d6a: char_row_bitmap <= 16'b1111111100000000;
		15'h4d6b: char_row_bitmap <= 16'b1111111100000000;
		15'h4d6c: char_row_bitmap <= 16'b1111111111111111;
		15'h4d6d: char_row_bitmap <= 16'b1111111111111111;
		15'h4d6e: char_row_bitmap <= 16'b1111111111111111;
		15'h4d6f: char_row_bitmap <= 16'b1111111111111111;
		15'h4d70: char_row_bitmap <= 16'b1111111111111111;
		15'h4d71: char_row_bitmap <= 16'b1111111111111111;
		15'h4d72: char_row_bitmap <= 16'b1111111111111111;
		15'h4d73: char_row_bitmap <= 16'b1111111111111111;
		15'h4d74: char_row_bitmap <= 16'b1111111111111111;
		15'h4d75: char_row_bitmap <= 16'b1111111111111111;
		15'h4d76: char_row_bitmap <= 16'b1111111111111111;
		15'h4d77: char_row_bitmap <= 16'b1111111111111111;
		15'h4d78: char_row_bitmap <= 16'b1111111111111111;
		15'h4d79: char_row_bitmap <= 16'b1111111111111111;
		15'h4d7a: char_row_bitmap <= 16'b1111111100000000;
		15'h4d7b: char_row_bitmap <= 16'b1111111100000000;
		15'h4d7c: char_row_bitmap <= 16'b1111111100000000;
		15'h4d7d: char_row_bitmap <= 16'b1111111100000000;
		15'h4d7e: char_row_bitmap <= 16'b1111111100000000;
		15'h4d7f: char_row_bitmap <= 16'b1111111100000000;
		15'h4d80: char_row_bitmap <= 16'b0000000000000000;
		15'h4d81: char_row_bitmap <= 16'b0000000000000000;
		15'h4d82: char_row_bitmap <= 16'b0000000000000000;
		15'h4d83: char_row_bitmap <= 16'b0000000000000000;
		15'h4d84: char_row_bitmap <= 16'b0000000000000000;
		15'h4d85: char_row_bitmap <= 16'b0000000000000000;
		15'h4d86: char_row_bitmap <= 16'b0000000000000000;
		15'h4d87: char_row_bitmap <= 16'b0000000000000000;
		15'h4d88: char_row_bitmap <= 16'b0000000000000000;
		15'h4d89: char_row_bitmap <= 16'b0000000000000000;
		15'h4d8a: char_row_bitmap <= 16'b0000000000000000;
		15'h4d8b: char_row_bitmap <= 16'b0000000000000000;
		15'h4d8c: char_row_bitmap <= 16'b0000000000000000;
		15'h4d8d: char_row_bitmap <= 16'b0000000000000000;
		15'h4d8e: char_row_bitmap <= 16'b0000000011111111;
		15'h4d8f: char_row_bitmap <= 16'b0000000011111111;
		15'h4d90: char_row_bitmap <= 16'b0000000011111111;
		15'h4d91: char_row_bitmap <= 16'b0000000011111111;
		15'h4d92: char_row_bitmap <= 16'b0000000011111111;
		15'h4d93: char_row_bitmap <= 16'b0000000011111111;
		15'h4d94: char_row_bitmap <= 16'b1111111100000000;
		15'h4d95: char_row_bitmap <= 16'b1111111100000000;
		15'h4d96: char_row_bitmap <= 16'b1111111100000000;
		15'h4d97: char_row_bitmap <= 16'b1111111100000000;
		15'h4d98: char_row_bitmap <= 16'b1111111100000000;
		15'h4d99: char_row_bitmap <= 16'b1111111100000000;
		15'h4d9a: char_row_bitmap <= 16'b0000000000000000;
		15'h4d9b: char_row_bitmap <= 16'b0000000000000000;
		15'h4d9c: char_row_bitmap <= 16'b0000000000000000;
		15'h4d9d: char_row_bitmap <= 16'b0000000000000000;
		15'h4d9e: char_row_bitmap <= 16'b0000000000000000;
		15'h4d9f: char_row_bitmap <= 16'b0000000000000000;
		15'h4da0: char_row_bitmap <= 16'b0000000000000000;
		15'h4da1: char_row_bitmap <= 16'b0000000000000000;
		15'h4da2: char_row_bitmap <= 16'b0000000011111111;
		15'h4da3: char_row_bitmap <= 16'b0000000011111111;
		15'h4da4: char_row_bitmap <= 16'b0000000011111111;
		15'h4da5: char_row_bitmap <= 16'b0000000011111111;
		15'h4da6: char_row_bitmap <= 16'b0000000011111111;
		15'h4da7: char_row_bitmap <= 16'b0000000011111111;
		15'h4da8: char_row_bitmap <= 16'b0000000011111111;
		15'h4da9: char_row_bitmap <= 16'b0000000011111111;
		15'h4daa: char_row_bitmap <= 16'b0000000011111111;
		15'h4dab: char_row_bitmap <= 16'b0000000011111111;
		15'h4dac: char_row_bitmap <= 16'b0000000011111111;
		15'h4dad: char_row_bitmap <= 16'b0000000011111111;
		15'h4dae: char_row_bitmap <= 16'b0000000000000000;
		15'h4daf: char_row_bitmap <= 16'b0000000000000000;
		15'h4db0: char_row_bitmap <= 16'b0000000000000000;
		15'h4db1: char_row_bitmap <= 16'b0000000000000000;
		15'h4db2: char_row_bitmap <= 16'b0000000000000000;
		15'h4db3: char_row_bitmap <= 16'b0000000000000000;
		15'h4db4: char_row_bitmap <= 16'b0000000000000000;
		15'h4db5: char_row_bitmap <= 16'b0000000000000000;
		15'h4db6: char_row_bitmap <= 16'b0000000011111111;
		15'h4db7: char_row_bitmap <= 16'b0000000011111111;
		15'h4db8: char_row_bitmap <= 16'b0000000011111111;
		15'h4db9: char_row_bitmap <= 16'b0000000011111111;
		15'h4dba: char_row_bitmap <= 16'b0000000011111111;
		15'h4dbb: char_row_bitmap <= 16'b0000000011111111;
		15'h4dbc: char_row_bitmap <= 16'b1111111111111111;
		15'h4dbd: char_row_bitmap <= 16'b1111111111111111;
		15'h4dbe: char_row_bitmap <= 16'b1111111111111111;
		15'h4dbf: char_row_bitmap <= 16'b1111111111111111;
		15'h4dc0: char_row_bitmap <= 16'b1111111111111111;
		15'h4dc1: char_row_bitmap <= 16'b1111111111111111;
		15'h4dc2: char_row_bitmap <= 16'b0000000000000000;
		15'h4dc3: char_row_bitmap <= 16'b0000000000000000;
		15'h4dc4: char_row_bitmap <= 16'b0000000000000000;
		15'h4dc5: char_row_bitmap <= 16'b0000000000000000;
		15'h4dc6: char_row_bitmap <= 16'b0000000000000000;
		15'h4dc7: char_row_bitmap <= 16'b0000000000000000;
		15'h4dc8: char_row_bitmap <= 16'b0000000000000000;
		15'h4dc9: char_row_bitmap <= 16'b0000000000000000;
		15'h4dca: char_row_bitmap <= 16'b0000000011111111;
		15'h4dcb: char_row_bitmap <= 16'b0000000011111111;
		15'h4dcc: char_row_bitmap <= 16'b0000000011111111;
		15'h4dcd: char_row_bitmap <= 16'b0000000011111111;
		15'h4dce: char_row_bitmap <= 16'b0000000011111111;
		15'h4dcf: char_row_bitmap <= 16'b0000000011111111;
		15'h4dd0: char_row_bitmap <= 16'b0000000000000000;
		15'h4dd1: char_row_bitmap <= 16'b0000000000000000;
		15'h4dd2: char_row_bitmap <= 16'b0000000000000000;
		15'h4dd3: char_row_bitmap <= 16'b0000000000000000;
		15'h4dd4: char_row_bitmap <= 16'b0000000000000000;
		15'h4dd5: char_row_bitmap <= 16'b0000000000000000;
		15'h4dd6: char_row_bitmap <= 16'b1111111100000000;
		15'h4dd7: char_row_bitmap <= 16'b1111111100000000;
		15'h4dd8: char_row_bitmap <= 16'b1111111100000000;
		15'h4dd9: char_row_bitmap <= 16'b1111111100000000;
		15'h4dda: char_row_bitmap <= 16'b1111111100000000;
		15'h4ddb: char_row_bitmap <= 16'b1111111100000000;
		15'h4ddc: char_row_bitmap <= 16'b1111111100000000;
		15'h4ddd: char_row_bitmap <= 16'b1111111100000000;
		15'h4dde: char_row_bitmap <= 16'b0000000011111111;
		15'h4ddf: char_row_bitmap <= 16'b0000000011111111;
		15'h4de0: char_row_bitmap <= 16'b0000000011111111;
		15'h4de1: char_row_bitmap <= 16'b0000000011111111;
		15'h4de2: char_row_bitmap <= 16'b0000000011111111;
		15'h4de3: char_row_bitmap <= 16'b0000000011111111;
		15'h4de4: char_row_bitmap <= 16'b1111111100000000;
		15'h4de5: char_row_bitmap <= 16'b1111111100000000;
		15'h4de6: char_row_bitmap <= 16'b1111111100000000;
		15'h4de7: char_row_bitmap <= 16'b1111111100000000;
		15'h4de8: char_row_bitmap <= 16'b1111111100000000;
		15'h4de9: char_row_bitmap <= 16'b1111111100000000;
		15'h4dea: char_row_bitmap <= 16'b1111111100000000;
		15'h4deb: char_row_bitmap <= 16'b1111111100000000;
		15'h4dec: char_row_bitmap <= 16'b1111111100000000;
		15'h4ded: char_row_bitmap <= 16'b1111111100000000;
		15'h4dee: char_row_bitmap <= 16'b1111111100000000;
		15'h4def: char_row_bitmap <= 16'b1111111100000000;
		15'h4df0: char_row_bitmap <= 16'b1111111100000000;
		15'h4df1: char_row_bitmap <= 16'b1111111100000000;
		15'h4df2: char_row_bitmap <= 16'b0000000011111111;
		15'h4df3: char_row_bitmap <= 16'b0000000011111111;
		15'h4df4: char_row_bitmap <= 16'b0000000011111111;
		15'h4df5: char_row_bitmap <= 16'b0000000011111111;
		15'h4df6: char_row_bitmap <= 16'b0000000011111111;
		15'h4df7: char_row_bitmap <= 16'b0000000011111111;
		15'h4df8: char_row_bitmap <= 16'b0000000011111111;
		15'h4df9: char_row_bitmap <= 16'b0000000011111111;
		15'h4dfa: char_row_bitmap <= 16'b0000000011111111;
		15'h4dfb: char_row_bitmap <= 16'b0000000011111111;
		15'h4dfc: char_row_bitmap <= 16'b0000000011111111;
		15'h4dfd: char_row_bitmap <= 16'b0000000011111111;
		15'h4dfe: char_row_bitmap <= 16'b1111111100000000;
		15'h4dff: char_row_bitmap <= 16'b1111111100000000;
		15'h4e00: char_row_bitmap <= 16'b1111111100000000;
		15'h4e01: char_row_bitmap <= 16'b1111111100000000;
		15'h4e02: char_row_bitmap <= 16'b1111111100000000;
		15'h4e03: char_row_bitmap <= 16'b1111111100000000;
		15'h4e04: char_row_bitmap <= 16'b1111111100000000;
		15'h4e05: char_row_bitmap <= 16'b1111111100000000;
		15'h4e06: char_row_bitmap <= 16'b0000000011111111;
		15'h4e07: char_row_bitmap <= 16'b0000000011111111;
		15'h4e08: char_row_bitmap <= 16'b0000000011111111;
		15'h4e09: char_row_bitmap <= 16'b0000000011111111;
		15'h4e0a: char_row_bitmap <= 16'b0000000011111111;
		15'h4e0b: char_row_bitmap <= 16'b0000000011111111;
		15'h4e0c: char_row_bitmap <= 16'b1111111111111111;
		15'h4e0d: char_row_bitmap <= 16'b1111111111111111;
		15'h4e0e: char_row_bitmap <= 16'b1111111111111111;
		15'h4e0f: char_row_bitmap <= 16'b1111111111111111;
		15'h4e10: char_row_bitmap <= 16'b1111111111111111;
		15'h4e11: char_row_bitmap <= 16'b1111111111111111;
		15'h4e12: char_row_bitmap <= 16'b1111111100000000;
		15'h4e13: char_row_bitmap <= 16'b1111111100000000;
		15'h4e14: char_row_bitmap <= 16'b1111111100000000;
		15'h4e15: char_row_bitmap <= 16'b1111111100000000;
		15'h4e16: char_row_bitmap <= 16'b1111111100000000;
		15'h4e17: char_row_bitmap <= 16'b1111111100000000;
		15'h4e18: char_row_bitmap <= 16'b1111111100000000;
		15'h4e19: char_row_bitmap <= 16'b1111111100000000;
		15'h4e1a: char_row_bitmap <= 16'b0000000011111111;
		15'h4e1b: char_row_bitmap <= 16'b0000000011111111;
		15'h4e1c: char_row_bitmap <= 16'b0000000011111111;
		15'h4e1d: char_row_bitmap <= 16'b0000000011111111;
		15'h4e1e: char_row_bitmap <= 16'b0000000011111111;
		15'h4e1f: char_row_bitmap <= 16'b0000000011111111;
		15'h4e20: char_row_bitmap <= 16'b0000000000000000;
		15'h4e21: char_row_bitmap <= 16'b0000000000000000;
		15'h4e22: char_row_bitmap <= 16'b0000000000000000;
		15'h4e23: char_row_bitmap <= 16'b0000000000000000;
		15'h4e24: char_row_bitmap <= 16'b0000000000000000;
		15'h4e25: char_row_bitmap <= 16'b0000000000000000;
		15'h4e26: char_row_bitmap <= 16'b0000000011111111;
		15'h4e27: char_row_bitmap <= 16'b0000000011111111;
		15'h4e28: char_row_bitmap <= 16'b0000000011111111;
		15'h4e29: char_row_bitmap <= 16'b0000000011111111;
		15'h4e2a: char_row_bitmap <= 16'b0000000011111111;
		15'h4e2b: char_row_bitmap <= 16'b0000000011111111;
		15'h4e2c: char_row_bitmap <= 16'b0000000011111111;
		15'h4e2d: char_row_bitmap <= 16'b0000000011111111;
		15'h4e2e: char_row_bitmap <= 16'b0000000011111111;
		15'h4e2f: char_row_bitmap <= 16'b0000000011111111;
		15'h4e30: char_row_bitmap <= 16'b0000000011111111;
		15'h4e31: char_row_bitmap <= 16'b0000000011111111;
		15'h4e32: char_row_bitmap <= 16'b0000000011111111;
		15'h4e33: char_row_bitmap <= 16'b0000000011111111;
		15'h4e34: char_row_bitmap <= 16'b1111111100000000;
		15'h4e35: char_row_bitmap <= 16'b1111111100000000;
		15'h4e36: char_row_bitmap <= 16'b1111111100000000;
		15'h4e37: char_row_bitmap <= 16'b1111111100000000;
		15'h4e38: char_row_bitmap <= 16'b1111111100000000;
		15'h4e39: char_row_bitmap <= 16'b1111111100000000;
		15'h4e3a: char_row_bitmap <= 16'b0000000011111111;
		15'h4e3b: char_row_bitmap <= 16'b0000000011111111;
		15'h4e3c: char_row_bitmap <= 16'b0000000011111111;
		15'h4e3d: char_row_bitmap <= 16'b0000000011111111;
		15'h4e3e: char_row_bitmap <= 16'b0000000011111111;
		15'h4e3f: char_row_bitmap <= 16'b0000000011111111;
		15'h4e40: char_row_bitmap <= 16'b0000000011111111;
		15'h4e41: char_row_bitmap <= 16'b0000000011111111;
		15'h4e42: char_row_bitmap <= 16'b0000000011111111;
		15'h4e43: char_row_bitmap <= 16'b0000000011111111;
		15'h4e44: char_row_bitmap <= 16'b0000000011111111;
		15'h4e45: char_row_bitmap <= 16'b0000000011111111;
		15'h4e46: char_row_bitmap <= 16'b0000000011111111;
		15'h4e47: char_row_bitmap <= 16'b0000000011111111;
		15'h4e48: char_row_bitmap <= 16'b0000000011111111;
		15'h4e49: char_row_bitmap <= 16'b0000000011111111;
		15'h4e4a: char_row_bitmap <= 16'b0000000011111111;
		15'h4e4b: char_row_bitmap <= 16'b0000000011111111;
		15'h4e4c: char_row_bitmap <= 16'b0000000011111111;
		15'h4e4d: char_row_bitmap <= 16'b0000000011111111;
		15'h4e4e: char_row_bitmap <= 16'b0000000011111111;
		15'h4e4f: char_row_bitmap <= 16'b0000000011111111;
		15'h4e50: char_row_bitmap <= 16'b0000000011111111;
		15'h4e51: char_row_bitmap <= 16'b0000000011111111;
		15'h4e52: char_row_bitmap <= 16'b0000000011111111;
		15'h4e53: char_row_bitmap <= 16'b0000000011111111;
		15'h4e54: char_row_bitmap <= 16'b0000000011111111;
		15'h4e55: char_row_bitmap <= 16'b0000000011111111;
		15'h4e56: char_row_bitmap <= 16'b0000000011111111;
		15'h4e57: char_row_bitmap <= 16'b0000000011111111;
		15'h4e58: char_row_bitmap <= 16'b0000000011111111;
		15'h4e59: char_row_bitmap <= 16'b0000000011111111;
		15'h4e5a: char_row_bitmap <= 16'b0000000011111111;
		15'h4e5b: char_row_bitmap <= 16'b0000000011111111;
		15'h4e5c: char_row_bitmap <= 16'b1111111111111111;
		15'h4e5d: char_row_bitmap <= 16'b1111111111111111;
		15'h4e5e: char_row_bitmap <= 16'b1111111111111111;
		15'h4e5f: char_row_bitmap <= 16'b1111111111111111;
		15'h4e60: char_row_bitmap <= 16'b1111111111111111;
		15'h4e61: char_row_bitmap <= 16'b1111111111111111;
		15'h4e62: char_row_bitmap <= 16'b0000000011111111;
		15'h4e63: char_row_bitmap <= 16'b0000000011111111;
		15'h4e64: char_row_bitmap <= 16'b0000000011111111;
		15'h4e65: char_row_bitmap <= 16'b0000000011111111;
		15'h4e66: char_row_bitmap <= 16'b0000000011111111;
		15'h4e67: char_row_bitmap <= 16'b0000000011111111;
		15'h4e68: char_row_bitmap <= 16'b0000000011111111;
		15'h4e69: char_row_bitmap <= 16'b0000000011111111;
		15'h4e6a: char_row_bitmap <= 16'b0000000011111111;
		15'h4e6b: char_row_bitmap <= 16'b0000000011111111;
		15'h4e6c: char_row_bitmap <= 16'b0000000011111111;
		15'h4e6d: char_row_bitmap <= 16'b0000000011111111;
		15'h4e6e: char_row_bitmap <= 16'b0000000011111111;
		15'h4e6f: char_row_bitmap <= 16'b0000000011111111;
		15'h4e70: char_row_bitmap <= 16'b0000000000000000;
		15'h4e71: char_row_bitmap <= 16'b0000000000000000;
		15'h4e72: char_row_bitmap <= 16'b0000000000000000;
		15'h4e73: char_row_bitmap <= 16'b0000000000000000;
		15'h4e74: char_row_bitmap <= 16'b0000000000000000;
		15'h4e75: char_row_bitmap <= 16'b0000000000000000;
		15'h4e76: char_row_bitmap <= 16'b1111111111111111;
		15'h4e77: char_row_bitmap <= 16'b1111111111111111;
		15'h4e78: char_row_bitmap <= 16'b1111111111111111;
		15'h4e79: char_row_bitmap <= 16'b1111111111111111;
		15'h4e7a: char_row_bitmap <= 16'b1111111111111111;
		15'h4e7b: char_row_bitmap <= 16'b1111111111111111;
		15'h4e7c: char_row_bitmap <= 16'b1111111111111111;
		15'h4e7d: char_row_bitmap <= 16'b1111111111111111;
		15'h4e7e: char_row_bitmap <= 16'b0000000011111111;
		15'h4e7f: char_row_bitmap <= 16'b0000000011111111;
		15'h4e80: char_row_bitmap <= 16'b0000000011111111;
		15'h4e81: char_row_bitmap <= 16'b0000000011111111;
		15'h4e82: char_row_bitmap <= 16'b0000000011111111;
		15'h4e83: char_row_bitmap <= 16'b0000000011111111;
		15'h4e84: char_row_bitmap <= 16'b1111111100000000;
		15'h4e85: char_row_bitmap <= 16'b1111111100000000;
		15'h4e86: char_row_bitmap <= 16'b1111111100000000;
		15'h4e87: char_row_bitmap <= 16'b1111111100000000;
		15'h4e88: char_row_bitmap <= 16'b1111111100000000;
		15'h4e89: char_row_bitmap <= 16'b1111111100000000;
		15'h4e8a: char_row_bitmap <= 16'b1111111111111111;
		15'h4e8b: char_row_bitmap <= 16'b1111111111111111;
		15'h4e8c: char_row_bitmap <= 16'b1111111111111111;
		15'h4e8d: char_row_bitmap <= 16'b1111111111111111;
		15'h4e8e: char_row_bitmap <= 16'b1111111111111111;
		15'h4e8f: char_row_bitmap <= 16'b1111111111111111;
		15'h4e90: char_row_bitmap <= 16'b1111111111111111;
		15'h4e91: char_row_bitmap <= 16'b1111111111111111;
		15'h4e92: char_row_bitmap <= 16'b0000000011111111;
		15'h4e93: char_row_bitmap <= 16'b0000000011111111;
		15'h4e94: char_row_bitmap <= 16'b0000000011111111;
		15'h4e95: char_row_bitmap <= 16'b0000000011111111;
		15'h4e96: char_row_bitmap <= 16'b0000000011111111;
		15'h4e97: char_row_bitmap <= 16'b0000000011111111;
		15'h4e98: char_row_bitmap <= 16'b0000000011111111;
		15'h4e99: char_row_bitmap <= 16'b0000000011111111;
		15'h4e9a: char_row_bitmap <= 16'b0000000011111111;
		15'h4e9b: char_row_bitmap <= 16'b0000000011111111;
		15'h4e9c: char_row_bitmap <= 16'b0000000011111111;
		15'h4e9d: char_row_bitmap <= 16'b0000000011111111;
		15'h4e9e: char_row_bitmap <= 16'b1111111111111111;
		15'h4e9f: char_row_bitmap <= 16'b1111111111111111;
		15'h4ea0: char_row_bitmap <= 16'b1111111111111111;
		15'h4ea1: char_row_bitmap <= 16'b1111111111111111;
		15'h4ea2: char_row_bitmap <= 16'b1111111111111111;
		15'h4ea3: char_row_bitmap <= 16'b1111111111111111;
		15'h4ea4: char_row_bitmap <= 16'b1111111111111111;
		15'h4ea5: char_row_bitmap <= 16'b1111111111111111;
		15'h4ea6: char_row_bitmap <= 16'b0000000011111111;
		15'h4ea7: char_row_bitmap <= 16'b0000000011111111;
		15'h4ea8: char_row_bitmap <= 16'b0000000011111111;
		15'h4ea9: char_row_bitmap <= 16'b0000000011111111;
		15'h4eaa: char_row_bitmap <= 16'b0000000011111111;
		15'h4eab: char_row_bitmap <= 16'b0000000011111111;
		15'h4eac: char_row_bitmap <= 16'b1111111111111111;
		15'h4ead: char_row_bitmap <= 16'b1111111111111111;
		15'h4eae: char_row_bitmap <= 16'b1111111111111111;
		15'h4eaf: char_row_bitmap <= 16'b1111111111111111;
		15'h4eb0: char_row_bitmap <= 16'b1111111111111111;
		15'h4eb1: char_row_bitmap <= 16'b1111111111111111;
		15'h4eb2: char_row_bitmap <= 16'b1111111111111111;
		15'h4eb3: char_row_bitmap <= 16'b1111111111111111;
		15'h4eb4: char_row_bitmap <= 16'b1111111111111111;
		15'h4eb5: char_row_bitmap <= 16'b1111111111111111;
		15'h4eb6: char_row_bitmap <= 16'b1111111111111111;
		15'h4eb7: char_row_bitmap <= 16'b1111111111111111;
		15'h4eb8: char_row_bitmap <= 16'b1111111111111111;
		15'h4eb9: char_row_bitmap <= 16'b1111111111111111;
		15'h4eba: char_row_bitmap <= 16'b0000000011111111;
		15'h4ebb: char_row_bitmap <= 16'b0000000011111111;
		15'h4ebc: char_row_bitmap <= 16'b0000000011111111;
		15'h4ebd: char_row_bitmap <= 16'b0000000011111111;
		15'h4ebe: char_row_bitmap <= 16'b0000000011111111;
		15'h4ebf: char_row_bitmap <= 16'b0000000011111111;
		15'h4ec0: char_row_bitmap <= 16'b0000000000000000;
		15'h4ec1: char_row_bitmap <= 16'b0000000000000000;
		15'h4ec2: char_row_bitmap <= 16'b0000000000000000;
		15'h4ec3: char_row_bitmap <= 16'b0000000000000000;
		15'h4ec4: char_row_bitmap <= 16'b0000000000000000;
		15'h4ec5: char_row_bitmap <= 16'b0000000000000000;
		15'h4ec6: char_row_bitmap <= 16'b0000000000000000;
		15'h4ec7: char_row_bitmap <= 16'b0000000000000000;
		15'h4ec8: char_row_bitmap <= 16'b0000000000000000;
		15'h4ec9: char_row_bitmap <= 16'b0000000000000000;
		15'h4eca: char_row_bitmap <= 16'b0000000000000000;
		15'h4ecb: char_row_bitmap <= 16'b0000000000000000;
		15'h4ecc: char_row_bitmap <= 16'b0000000000000000;
		15'h4ecd: char_row_bitmap <= 16'b0000000000000000;
		15'h4ece: char_row_bitmap <= 16'b1111111111111111;
		15'h4ecf: char_row_bitmap <= 16'b1111111111111111;
		15'h4ed0: char_row_bitmap <= 16'b1111111111111111;
		15'h4ed1: char_row_bitmap <= 16'b1111111111111111;
		15'h4ed2: char_row_bitmap <= 16'b1111111111111111;
		15'h4ed3: char_row_bitmap <= 16'b1111111111111111;
		15'h4ed4: char_row_bitmap <= 16'b1111111100000000;
		15'h4ed5: char_row_bitmap <= 16'b1111111100000000;
		15'h4ed6: char_row_bitmap <= 16'b1111111100000000;
		15'h4ed7: char_row_bitmap <= 16'b1111111100000000;
		15'h4ed8: char_row_bitmap <= 16'b1111111100000000;
		15'h4ed9: char_row_bitmap <= 16'b1111111100000000;
		15'h4eda: char_row_bitmap <= 16'b0000000000000000;
		15'h4edb: char_row_bitmap <= 16'b0000000000000000;
		15'h4edc: char_row_bitmap <= 16'b0000000000000000;
		15'h4edd: char_row_bitmap <= 16'b0000000000000000;
		15'h4ede: char_row_bitmap <= 16'b0000000000000000;
		15'h4edf: char_row_bitmap <= 16'b0000000000000000;
		15'h4ee0: char_row_bitmap <= 16'b0000000000000000;
		15'h4ee1: char_row_bitmap <= 16'b0000000000000000;
		15'h4ee2: char_row_bitmap <= 16'b1111111111111111;
		15'h4ee3: char_row_bitmap <= 16'b1111111111111111;
		15'h4ee4: char_row_bitmap <= 16'b1111111111111111;
		15'h4ee5: char_row_bitmap <= 16'b1111111111111111;
		15'h4ee6: char_row_bitmap <= 16'b1111111111111111;
		15'h4ee7: char_row_bitmap <= 16'b1111111111111111;
		15'h4ee8: char_row_bitmap <= 16'b0000000011111111;
		15'h4ee9: char_row_bitmap <= 16'b0000000011111111;
		15'h4eea: char_row_bitmap <= 16'b0000000011111111;
		15'h4eeb: char_row_bitmap <= 16'b0000000011111111;
		15'h4eec: char_row_bitmap <= 16'b0000000011111111;
		15'h4eed: char_row_bitmap <= 16'b0000000011111111;
		15'h4eee: char_row_bitmap <= 16'b0000000000000000;
		15'h4eef: char_row_bitmap <= 16'b0000000000000000;
		15'h4ef0: char_row_bitmap <= 16'b0000000000000000;
		15'h4ef1: char_row_bitmap <= 16'b0000000000000000;
		15'h4ef2: char_row_bitmap <= 16'b0000000000000000;
		15'h4ef3: char_row_bitmap <= 16'b0000000000000000;
		15'h4ef4: char_row_bitmap <= 16'b0000000000000000;
		15'h4ef5: char_row_bitmap <= 16'b0000000000000000;
		15'h4ef6: char_row_bitmap <= 16'b1111111111111111;
		15'h4ef7: char_row_bitmap <= 16'b1111111111111111;
		15'h4ef8: char_row_bitmap <= 16'b1111111111111111;
		15'h4ef9: char_row_bitmap <= 16'b1111111111111111;
		15'h4efa: char_row_bitmap <= 16'b1111111111111111;
		15'h4efb: char_row_bitmap <= 16'b1111111111111111;
		15'h4efc: char_row_bitmap <= 16'b1111111111111111;
		15'h4efd: char_row_bitmap <= 16'b1111111111111111;
		15'h4efe: char_row_bitmap <= 16'b1111111111111111;
		15'h4eff: char_row_bitmap <= 16'b1111111111111111;
		15'h4f00: char_row_bitmap <= 16'b1111111111111111;
		15'h4f01: char_row_bitmap <= 16'b1111111111111111;
		15'h4f02: char_row_bitmap <= 16'b0000000000000000;
		15'h4f03: char_row_bitmap <= 16'b0000000000000000;
		15'h4f04: char_row_bitmap <= 16'b0000000000000000;
		15'h4f05: char_row_bitmap <= 16'b0000000000000000;
		15'h4f06: char_row_bitmap <= 16'b0000000000000000;
		15'h4f07: char_row_bitmap <= 16'b0000000000000000;
		15'h4f08: char_row_bitmap <= 16'b0000000000000000;
		15'h4f09: char_row_bitmap <= 16'b0000000000000000;
		15'h4f0a: char_row_bitmap <= 16'b1111111111111111;
		15'h4f0b: char_row_bitmap <= 16'b1111111111111111;
		15'h4f0c: char_row_bitmap <= 16'b1111111111111111;
		15'h4f0d: char_row_bitmap <= 16'b1111111111111111;
		15'h4f0e: char_row_bitmap <= 16'b1111111111111111;
		15'h4f0f: char_row_bitmap <= 16'b1111111111111111;
		15'h4f10: char_row_bitmap <= 16'b0000000000000000;
		15'h4f11: char_row_bitmap <= 16'b0000000000000000;
		15'h4f12: char_row_bitmap <= 16'b0000000000000000;
		15'h4f13: char_row_bitmap <= 16'b0000000000000000;
		15'h4f14: char_row_bitmap <= 16'b0000000000000000;
		15'h4f15: char_row_bitmap <= 16'b0000000000000000;
		15'h4f16: char_row_bitmap <= 16'b1111111100000000;
		15'h4f17: char_row_bitmap <= 16'b1111111100000000;
		15'h4f18: char_row_bitmap <= 16'b1111111100000000;
		15'h4f19: char_row_bitmap <= 16'b1111111100000000;
		15'h4f1a: char_row_bitmap <= 16'b1111111100000000;
		15'h4f1b: char_row_bitmap <= 16'b1111111100000000;
		15'h4f1c: char_row_bitmap <= 16'b1111111100000000;
		15'h4f1d: char_row_bitmap <= 16'b1111111100000000;
		15'h4f1e: char_row_bitmap <= 16'b1111111111111111;
		15'h4f1f: char_row_bitmap <= 16'b1111111111111111;
		15'h4f20: char_row_bitmap <= 16'b1111111111111111;
		15'h4f21: char_row_bitmap <= 16'b1111111111111111;
		15'h4f22: char_row_bitmap <= 16'b1111111111111111;
		15'h4f23: char_row_bitmap <= 16'b1111111111111111;
		15'h4f24: char_row_bitmap <= 16'b1111111100000000;
		15'h4f25: char_row_bitmap <= 16'b1111111100000000;
		15'h4f26: char_row_bitmap <= 16'b1111111100000000;
		15'h4f27: char_row_bitmap <= 16'b1111111100000000;
		15'h4f28: char_row_bitmap <= 16'b1111111100000000;
		15'h4f29: char_row_bitmap <= 16'b1111111100000000;
		15'h4f2a: char_row_bitmap <= 16'b1111111100000000;
		15'h4f2b: char_row_bitmap <= 16'b1111111100000000;
		15'h4f2c: char_row_bitmap <= 16'b1111111100000000;
		15'h4f2d: char_row_bitmap <= 16'b1111111100000000;
		15'h4f2e: char_row_bitmap <= 16'b1111111100000000;
		15'h4f2f: char_row_bitmap <= 16'b1111111100000000;
		15'h4f30: char_row_bitmap <= 16'b1111111100000000;
		15'h4f31: char_row_bitmap <= 16'b1111111100000000;
		15'h4f32: char_row_bitmap <= 16'b1111111111111111;
		15'h4f33: char_row_bitmap <= 16'b1111111111111111;
		15'h4f34: char_row_bitmap <= 16'b1111111111111111;
		15'h4f35: char_row_bitmap <= 16'b1111111111111111;
		15'h4f36: char_row_bitmap <= 16'b1111111111111111;
		15'h4f37: char_row_bitmap <= 16'b1111111111111111;
		15'h4f38: char_row_bitmap <= 16'b0000000011111111;
		15'h4f39: char_row_bitmap <= 16'b0000000011111111;
		15'h4f3a: char_row_bitmap <= 16'b0000000011111111;
		15'h4f3b: char_row_bitmap <= 16'b0000000011111111;
		15'h4f3c: char_row_bitmap <= 16'b0000000011111111;
		15'h4f3d: char_row_bitmap <= 16'b0000000011111111;
		15'h4f3e: char_row_bitmap <= 16'b1111111100000000;
		15'h4f3f: char_row_bitmap <= 16'b1111111100000000;
		15'h4f40: char_row_bitmap <= 16'b1111111100000000;
		15'h4f41: char_row_bitmap <= 16'b1111111100000000;
		15'h4f42: char_row_bitmap <= 16'b1111111100000000;
		15'h4f43: char_row_bitmap <= 16'b1111111100000000;
		15'h4f44: char_row_bitmap <= 16'b1111111100000000;
		15'h4f45: char_row_bitmap <= 16'b1111111100000000;
		15'h4f46: char_row_bitmap <= 16'b1111111111111111;
		15'h4f47: char_row_bitmap <= 16'b1111111111111111;
		15'h4f48: char_row_bitmap <= 16'b1111111111111111;
		15'h4f49: char_row_bitmap <= 16'b1111111111111111;
		15'h4f4a: char_row_bitmap <= 16'b1111111111111111;
		15'h4f4b: char_row_bitmap <= 16'b1111111111111111;
		15'h4f4c: char_row_bitmap <= 16'b1111111111111111;
		15'h4f4d: char_row_bitmap <= 16'b1111111111111111;
		15'h4f4e: char_row_bitmap <= 16'b1111111111111111;
		15'h4f4f: char_row_bitmap <= 16'b1111111111111111;
		15'h4f50: char_row_bitmap <= 16'b1111111111111111;
		15'h4f51: char_row_bitmap <= 16'b1111111111111111;
		15'h4f52: char_row_bitmap <= 16'b1111111100000000;
		15'h4f53: char_row_bitmap <= 16'b1111111100000000;
		15'h4f54: char_row_bitmap <= 16'b1111111100000000;
		15'h4f55: char_row_bitmap <= 16'b1111111100000000;
		15'h4f56: char_row_bitmap <= 16'b1111111100000000;
		15'h4f57: char_row_bitmap <= 16'b1111111100000000;
		15'h4f58: char_row_bitmap <= 16'b1111111100000000;
		15'h4f59: char_row_bitmap <= 16'b1111111100000000;
		15'h4f5a: char_row_bitmap <= 16'b1111111111111111;
		15'h4f5b: char_row_bitmap <= 16'b1111111111111111;
		15'h4f5c: char_row_bitmap <= 16'b1111111111111111;
		15'h4f5d: char_row_bitmap <= 16'b1111111111111111;
		15'h4f5e: char_row_bitmap <= 16'b1111111111111111;
		15'h4f5f: char_row_bitmap <= 16'b1111111111111111;
		15'h4f60: char_row_bitmap <= 16'b0000000000000000;
		15'h4f61: char_row_bitmap <= 16'b0000000000000000;
		15'h4f62: char_row_bitmap <= 16'b0000000000000000;
		15'h4f63: char_row_bitmap <= 16'b0000000000000000;
		15'h4f64: char_row_bitmap <= 16'b0000000000000000;
		15'h4f65: char_row_bitmap <= 16'b0000000000000000;
		15'h4f66: char_row_bitmap <= 16'b0000000011111111;
		15'h4f67: char_row_bitmap <= 16'b0000000011111111;
		15'h4f68: char_row_bitmap <= 16'b0000000011111111;
		15'h4f69: char_row_bitmap <= 16'b0000000011111111;
		15'h4f6a: char_row_bitmap <= 16'b0000000011111111;
		15'h4f6b: char_row_bitmap <= 16'b0000000011111111;
		15'h4f6c: char_row_bitmap <= 16'b0000000011111111;
		15'h4f6d: char_row_bitmap <= 16'b0000000011111111;
		15'h4f6e: char_row_bitmap <= 16'b1111111111111111;
		15'h4f6f: char_row_bitmap <= 16'b1111111111111111;
		15'h4f70: char_row_bitmap <= 16'b1111111111111111;
		15'h4f71: char_row_bitmap <= 16'b1111111111111111;
		15'h4f72: char_row_bitmap <= 16'b1111111111111111;
		15'h4f73: char_row_bitmap <= 16'b1111111111111111;
		15'h4f74: char_row_bitmap <= 16'b1111111100000000;
		15'h4f75: char_row_bitmap <= 16'b1111111100000000;
		15'h4f76: char_row_bitmap <= 16'b1111111100000000;
		15'h4f77: char_row_bitmap <= 16'b1111111100000000;
		15'h4f78: char_row_bitmap <= 16'b1111111100000000;
		15'h4f79: char_row_bitmap <= 16'b1111111100000000;
		15'h4f7a: char_row_bitmap <= 16'b0000000011111111;
		15'h4f7b: char_row_bitmap <= 16'b0000000011111111;
		15'h4f7c: char_row_bitmap <= 16'b0000000011111111;
		15'h4f7d: char_row_bitmap <= 16'b0000000011111111;
		15'h4f7e: char_row_bitmap <= 16'b0000000011111111;
		15'h4f7f: char_row_bitmap <= 16'b0000000011111111;
		15'h4f80: char_row_bitmap <= 16'b0000000011111111;
		15'h4f81: char_row_bitmap <= 16'b0000000011111111;
		15'h4f82: char_row_bitmap <= 16'b1111111111111111;
		15'h4f83: char_row_bitmap <= 16'b1111111111111111;
		15'h4f84: char_row_bitmap <= 16'b1111111111111111;
		15'h4f85: char_row_bitmap <= 16'b1111111111111111;
		15'h4f86: char_row_bitmap <= 16'b1111111111111111;
		15'h4f87: char_row_bitmap <= 16'b1111111111111111;
		15'h4f88: char_row_bitmap <= 16'b0000000011111111;
		15'h4f89: char_row_bitmap <= 16'b0000000011111111;
		15'h4f8a: char_row_bitmap <= 16'b0000000011111111;
		15'h4f8b: char_row_bitmap <= 16'b0000000011111111;
		15'h4f8c: char_row_bitmap <= 16'b0000000011111111;
		15'h4f8d: char_row_bitmap <= 16'b0000000011111111;
		15'h4f8e: char_row_bitmap <= 16'b0000000011111111;
		15'h4f8f: char_row_bitmap <= 16'b0000000011111111;
		15'h4f90: char_row_bitmap <= 16'b0000000011111111;
		15'h4f91: char_row_bitmap <= 16'b0000000011111111;
		15'h4f92: char_row_bitmap <= 16'b0000000011111111;
		15'h4f93: char_row_bitmap <= 16'b0000000011111111;
		15'h4f94: char_row_bitmap <= 16'b0000000011111111;
		15'h4f95: char_row_bitmap <= 16'b0000000011111111;
		15'h4f96: char_row_bitmap <= 16'b1111111111111111;
		15'h4f97: char_row_bitmap <= 16'b1111111111111111;
		15'h4f98: char_row_bitmap <= 16'b1111111111111111;
		15'h4f99: char_row_bitmap <= 16'b1111111111111111;
		15'h4f9a: char_row_bitmap <= 16'b1111111111111111;
		15'h4f9b: char_row_bitmap <= 16'b1111111111111111;
		15'h4f9c: char_row_bitmap <= 16'b1111111111111111;
		15'h4f9d: char_row_bitmap <= 16'b1111111111111111;
		15'h4f9e: char_row_bitmap <= 16'b1111111111111111;
		15'h4f9f: char_row_bitmap <= 16'b1111111111111111;
		15'h4fa0: char_row_bitmap <= 16'b1111111111111111;
		15'h4fa1: char_row_bitmap <= 16'b1111111111111111;
		15'h4fa2: char_row_bitmap <= 16'b0000000011111111;
		15'h4fa3: char_row_bitmap <= 16'b0000000011111111;
		15'h4fa4: char_row_bitmap <= 16'b0000000011111111;
		15'h4fa5: char_row_bitmap <= 16'b0000000011111111;
		15'h4fa6: char_row_bitmap <= 16'b0000000011111111;
		15'h4fa7: char_row_bitmap <= 16'b0000000011111111;
		15'h4fa8: char_row_bitmap <= 16'b0000000011111111;
		15'h4fa9: char_row_bitmap <= 16'b0000000011111111;
		15'h4faa: char_row_bitmap <= 16'b1111111111111111;
		15'h4fab: char_row_bitmap <= 16'b1111111111111111;
		15'h4fac: char_row_bitmap <= 16'b1111111111111111;
		15'h4fad: char_row_bitmap <= 16'b1111111111111111;
		15'h4fae: char_row_bitmap <= 16'b1111111111111111;
		15'h4faf: char_row_bitmap <= 16'b1111111111111111;
		15'h4fb0: char_row_bitmap <= 16'b0000000000000000;
		15'h4fb1: char_row_bitmap <= 16'b0000000000000000;
		15'h4fb2: char_row_bitmap <= 16'b0000000000000000;
		15'h4fb3: char_row_bitmap <= 16'b0000000000000000;
		15'h4fb4: char_row_bitmap <= 16'b0000000000000000;
		15'h4fb5: char_row_bitmap <= 16'b0000000000000000;
		15'h4fb6: char_row_bitmap <= 16'b1111111111111111;
		15'h4fb7: char_row_bitmap <= 16'b1111111111111111;
		15'h4fb8: char_row_bitmap <= 16'b1111111111111111;
		15'h4fb9: char_row_bitmap <= 16'b1111111111111111;
		15'h4fba: char_row_bitmap <= 16'b1111111111111111;
		15'h4fbb: char_row_bitmap <= 16'b1111111111111111;
		15'h4fbc: char_row_bitmap <= 16'b1111111111111111;
		15'h4fbd: char_row_bitmap <= 16'b1111111111111111;
		15'h4fbe: char_row_bitmap <= 16'b1111111111111111;
		15'h4fbf: char_row_bitmap <= 16'b1111111111111111;
		15'h4fc0: char_row_bitmap <= 16'b1111111111111111;
		15'h4fc1: char_row_bitmap <= 16'b1111111111111111;
		15'h4fc2: char_row_bitmap <= 16'b1111111111111111;
		15'h4fc3: char_row_bitmap <= 16'b1111111111111111;
		15'h4fc4: char_row_bitmap <= 16'b1111111100000000;
		15'h4fc5: char_row_bitmap <= 16'b1111111100000000;
		15'h4fc6: char_row_bitmap <= 16'b1111111100000000;
		15'h4fc7: char_row_bitmap <= 16'b1111111100000000;
		15'h4fc8: char_row_bitmap <= 16'b1111111100000000;
		15'h4fc9: char_row_bitmap <= 16'b1111111100000000;
		15'h4fca: char_row_bitmap <= 16'b1111111111111111;
		15'h4fcb: char_row_bitmap <= 16'b1111111111111111;
		15'h4fcc: char_row_bitmap <= 16'b1111111111111111;
		15'h4fcd: char_row_bitmap <= 16'b1111111111111111;
		15'h4fce: char_row_bitmap <= 16'b1111111111111111;
		15'h4fcf: char_row_bitmap <= 16'b1111111111111111;
		15'h4fd0: char_row_bitmap <= 16'b1111111111111111;
		15'h4fd1: char_row_bitmap <= 16'b1111111111111111;
		15'h4fd2: char_row_bitmap <= 16'b1111111111111111;
		15'h4fd3: char_row_bitmap <= 16'b1111111111111111;
		15'h4fd4: char_row_bitmap <= 16'b1111111111111111;
		15'h4fd5: char_row_bitmap <= 16'b1111111111111111;
		15'h4fd6: char_row_bitmap <= 16'b1111111111111111;
		15'h4fd7: char_row_bitmap <= 16'b1111111111111111;
		15'h4fd8: char_row_bitmap <= 16'b0000000011111111;
		15'h4fd9: char_row_bitmap <= 16'b0000000011111111;
		15'h4fda: char_row_bitmap <= 16'b0000000011111111;
		15'h4fdb: char_row_bitmap <= 16'b0000000011111111;
		15'h4fdc: char_row_bitmap <= 16'b0000000011111111;
		15'h4fdd: char_row_bitmap <= 16'b0000000011111111;
		15'h4fde: char_row_bitmap <= 16'b1111111111111111;
		15'h4fdf: char_row_bitmap <= 16'b1111111111111111;
		15'h4fe0: char_row_bitmap <= 16'b1111111111111111;
		15'h4fe1: char_row_bitmap <= 16'b1111111111111111;
		15'h4fe2: char_row_bitmap <= 16'b1111111111111111;
		15'h4fe3: char_row_bitmap <= 16'b1111111111111111;
		15'h4fe4: char_row_bitmap <= 16'b1111111111111111;
		15'h4fe5: char_row_bitmap <= 16'b1111111111111111;
		15'h4fe6: char_row_bitmap <= 16'b1111111111111111;
		15'h4fe7: char_row_bitmap <= 16'b1111111111111111;
		15'h4fe8: char_row_bitmap <= 16'b1111111111111111;
		15'h4fe9: char_row_bitmap <= 16'b1111111111111111;
		15'h4fea: char_row_bitmap <= 16'b1111111111111111;
		15'h4feb: char_row_bitmap <= 16'b1111111111111111;
		15'h4fec: char_row_bitmap <= 16'b1111111111111111;
		15'h4fed: char_row_bitmap <= 16'b1111111111111111;
		15'h4fee: char_row_bitmap <= 16'b1111111111111111;
		15'h4fef: char_row_bitmap <= 16'b1111111111111111;
		15'h4ff0: char_row_bitmap <= 16'b1111111111111111;
		15'h4ff1: char_row_bitmap <= 16'b1111111111111111;
		15'h4ff2: char_row_bitmap <= 16'b1111111111111111;
		15'h4ff3: char_row_bitmap <= 16'b1111111111111111;
		15'h4ff4: char_row_bitmap <= 16'b1111111111111111;
		15'h4ff5: char_row_bitmap <= 16'b1111111111111111;
		15'h4ff6: char_row_bitmap <= 16'b1111111111111111;
		15'h4ff7: char_row_bitmap <= 16'b1111111111111111;
		15'h4ff8: char_row_bitmap <= 16'b1111111111111111;
		15'h4ff9: char_row_bitmap <= 16'b1111111111111111;
		15'h4ffa: char_row_bitmap <= 16'b1111111111111111;
		15'h4ffb: char_row_bitmap <= 16'b1111111111111111;
		15'h4ffc: char_row_bitmap <= 16'b1111111111111111;
		15'h4ffd: char_row_bitmap <= 16'b1111111111111111;
		15'h4ffe: char_row_bitmap <= 16'b1111111111111111;
		15'h4fff: char_row_bitmap <= 16'b1111111111111111;
    endcase

endmodule

localparam
	TS_CURSOR_NOP = 'd0,
	TS_CURSOR_SET = 'd1,
	TS_CURSOR_UP = 'd2,
	TS_CURSOR_DOWN = 'd3,
	TS_CURSOR_LEFT = 'd4,
	TS_CURSOR_RIGHT = 'd5,
	TS_CURSOR_NEXT_CHAR = 'd6,
	TS_CURSOR_LINE_FEED = 'd7;

localparam
	TS_ORIENTATION_RIGHT = 'd0,
	TS_ORIENTATION_LEFT  = 'd1,
	TS_ORIENTATION_DOWN  = 'd2,
	TS_ORIENTATION_UP    = 'd3;

// Verilog netlist created by TD v4.6.25304
// Mon May 31 15:09:41 2021

`timescale 1ns / 1ps
module cursor_ram  // al_ip/cursor_ram.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [8:0] addra;  // al_ip/cursor_ram.v(18)
  input clka;  // al_ip/cursor_ram.v(19)
  input rsta;  // al_ip/cursor_ram.v(20)
  output [15:0] doa;  // al_ip/cursor_ram.v(16)


  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=384;width=16;num_section=1;width_per_section=16;section_size=16;working_depth=512;working_width=18;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("0"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("18"),
    .DATA_WIDTH_B("18"),
    .INITP_00(256'h0555555555555550000005000000011511111110044000100400400000001000),
    .INITP_01(256'h0000011400000000040114004110400000555554010000011444444500000000),
    .INITP_02(256'h0000000000000500005000000000000000000005050000000000000000000500),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000075AB000075AC000075B0000075C000007500000076000000780000006000),
    .INIT_01(256'h600075AA5FFC75AA55B075AA55C075AA550075AA560075AA580075AA600075AA),
    .INIT_02(256'h1E000000750000007500000056006003560078035800760E5800750E600075FA),
    .INIT_03(256'h000001AC000001AC000001AC000001AC000001AC000001AC000001AC000000F0),
    .INIT_04(256'h55AB1DAA55AB75AA55AB75AA55AB75AA55AB75AA5DEB75AE5DEC1DAE673007AF),
    .INIT_05(256'h00000000000000000000000000000000000000007FFC07FF55AC07AA55AB1DAA),
    .INIT_06(256'h2A7F7E552A7F7E557FFF7FFF7FFC1FFF7FFC1FFF7FF007FF7FC001FF7E00003F),
    .INIT_07(256'h7E00003F7FC001FF7FF007FF7FFC1FFF7FFC1FFF7FFF7FFF2A7F7E552A7F7E55),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h2E00066A55001DAA55001DAA55001DAA55001DAA55001DAA55001DAA7FC07FFF),
    .INIT_0A(256'h560007A6580001AA600000EA0000003B0000000C00000037600000D538000155),
    .INIT_0B(256'h00000000000000007FC07FFF2B001A552B001A552B001A552D001C5535001D55),
    .INIT_0C(256'h5FAC1DFE58F0070E58C0010E5800000E5F0000FE5600003A5800000E60000003),
    .INIT_0D(256'h5600003A5F0000FE5800000E58C0010E58F0070E5FAC1DFE55AB75AA55AB75AA),
    .INIT_0E(256'h000000000000000000000000000000000000000000000000600000035800000E),
    .INIT_0F(256'h55AB1DAA55AB75AA55AB75AA55AB75AA55AB75AA5DEB75AE5DEC1DAE673006F3),
    .INIT_10(256'h00000000000000000000000000000000000000007FFC07FF55AC07AA55AB1DAA),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h1DAC75B007F01FC0000000036000000E6000000E6000000E6000000E00000003),
    .INIT_13(256'h00000000000000036000000E6000000E6000000E6000000E0000000307F01FC0),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h55AB75AA55AB75AA57FC1FFA5600003A5600003A5600003A5600003A7800000F),
    .INIT_16(256'h7800000F5600003A5600003A5600003A5600003A57FC1FFA55AB75AA55AB75AA),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("PDPW8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_384x16_sub_000000_000 (
    .addra({addra,4'b1111}),
    .addrb({addra,4'b1111}),
    .clka(clka),
    .clkb(clka),
    .dia(9'b000000000),
    .dib({open_n55,open_n56,7'b0000000}),
    .rsta(rsta),
    .rstb(rsta),
    .doa(doa[8:0]),
    .dob({open_n61,open_n62,doa[15:9]}));

endmodule 

